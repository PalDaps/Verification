`ifndef OVM_AHB_VC_PKG
`define OVM_AHB_VC_PKG

`include "ahb_if.sv"

package ovm_ahb_vc_pkg;

   import ovm_pkg::*;
  `include "ovm_macros.svh"

  `include "ovm_ahb_vc_class_files.sv"

endpackage

`endif