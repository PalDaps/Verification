  
  `include "ovm_spi_if_wrapper.sv"
  `include "ovm_spi_tran_item.sv"
  `include "ovm_spi_slave_driver.sv"
  `include "ovm_spi_slave_sequencer.sv"
  `include "ovm_spi_seq_lib.sv"
  `include "ovm_spi_monitor.sv"
  `include "ovm_spi_agent.sv"