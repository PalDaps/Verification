import `uvm_ovm_(pkg)::*;

`ifndef UNILANG_OVM
  import cdns_uvm_pkg::*;
`endif

package unilang;
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
0EmVapT+EPc9jukwqT4dot0PfPb7FiXKF5HO7oXVJtnT3/rGAIvlVaF5pw6Lw3Ez
fJ2JOWyjt+HEM4Zf8JQNtxpfp4q86C7PzN+tiZQ99TDZ5vk52ropbhnrc6QR7Poe
hLTCtMF2uvZklKhcWlX5pfeyap8Rwa1VCjOPRZqC88hJul5auYiYcA==
//pragma protect end_key_block
//pragma protect digest_block
FCezBCW5uI6z/c2HXWALqQvz3oc=
//pragma protect end_digest_block
//pragma protect data_block
vQJgnjZfS5hdXtD3hV1bon8a4aZpGvRZDum5/HRvLnIU2TaM8P/fjJHjFPo+FWML
LUWKPuHu7sHr9ahbCj9DcQdof8/K2Uxt+xt/f4E1SmqBWfHeNYGc/9W0savZu3eN
8Gy78ITvA1F4qxIHwBNT7GCn/8EoVxDUFwvZYjzSD2msE+jvG99nkHopHZoxa9wy
hsdEiFTxI5AoqWo7bq8VqxQn+q4II1ORfVq2HiqeCOcNhHuo1Jz/3jkdS27VMerV
JubzQ0AeHxV3/9SLQBSKR5HnTtf8UpNMqR9yj1pI5aP+NZ0wzykfF3hcICBVjrEh
lR9nbHLbeJEuKgKQ8YZyQwvHa/9j5KAkBf8VVBAnFzxyk0yI2RcC0ldY7+8lPH7U
Smor1vZtUOxrjDZGWdRZVKL1VMw/dFjlx5CgOW9EGYZZU+U8G9om72tV3sqEfLBC
Koq31I1TJnLrymu0nzRbPYDJcQyfiGXaqox510MW108APfTkJi9MO+qeyiJF1qs1
PpB5RyceQ8dFgnAn7yAbekG/ZaEGu66NvaBUC1ARD118ayCfltzaT9lcr2rKHQO/
nejBkCQ7rrX2KOxdqnD9fB/lnojWbb3Av0an91USNapRP69Ag2eEKRNFMPvYRGYx
14DwIuZNNB/4TGHBnAqhEWR12rtJcV/3+1sNszbvq+mHjyvUJVK7Y5DqhxBDlgc2
48962JIcggf/qVeX4XA2dsbJebVdKaYq9FnSOTC+HedDdq76YVtRayiMJyyVWkKK
CLetzEe0B6xJncn/cqxh/pwEQmMn9NBwk8LpPCoqen0/W1ALm+MV0sBVzMKgqF3N
kvn2gf+Fss3WRqQszw158AvlzBMOf9gUNrK031jEyPl9J8awosL6JTTxEVlX0zI5
NfZ0ZSF3+/ktMp6FMfjs6HKVNiftzQJ9XOsL/P4S5ldwx03XDAQcw81eG+p1mXG3
wfqyIpM7a3Zs+LbtOIUoG5BJc9Pp8GbxnRyx6uGxIEF3MMLMUiO4s1d7TvPuPFdB
vrh0yLA9kXoze5ykbrj8aVQhwV8DlZmfGZHSnGNKIpCj8urNmD8UmT1xGdaTiP0J
PLuk/CxGjCsq3M6Kee1vDipD9Zb1UvwTiD7cRlPFag0lxCKeqbBdOHV2adHLkQsL
UtN7CstVQxb20xDSNJ2SpCLGCEH/T4KQFG7rDO1u1+rJuJOysVNy6NRwj3aVrc/C
nK55igq7rckZ/GXRVDCqs9EAa1DZmqf7uF3pbuB9aMjs+r25MTfYXreIUp2IsGcp
kTgdGKlWMLdilVPwfedGexf214bo1GuF5EqAZO2F+as7zCm6wB6YGo4ij1ZCop0d
BfUfzaTHfM6ItorLbKRTvHaQ1p1rFm6qgUHIC9Io6RGK2EBRSi172kx7TMPRd/Fo
7Wk4hBzY+uoR3GAtodXtmiKoTq8anVgeYrP6FTChS9YVGvMwVer+pux5SUUQZXdA
hxFQ7fCJX7twP2mO19i9YhefDiZ/eQ8AvS6IY3aAT1zwnm3Km1axBpzbiaVXjPx5
1G4QFHNLptV5X+S6uohyZcFUiyteZKG/ybH3MmN2iubHsXdTX4k+XLmA9niT6gZq
edhgGCDKNWS4Dzn0Ce4J4VKC9dY6gGjgSJ/uReYcMRo8NkTO7oyWFmxo2ye6O3J0
+lOzTBvHqjMkY/mrG6Kkyhx4fv++qTJ346uvgRwtTIfe0VGs/ngtX+BZsJxTTsKC
S9XsRqzTsRoVhsT6I4bIm78onMoPVkPU2m6D23f0+zDtp3PsSprwcneYAuV9/dfT
3R7bm70aqGQTdsX1nDUNKMMSs6xvcgArU3qCtUhZcIbKqYjrTi+AC3hthLMr+V8Y
nLsouZMdCwDsjmS95OrBFDcY40GZBmzupwmgBIgOlK3wpELIhWNCa0sZuulKgEJx
RYyG+JsQxJ9J02hzNDLPShg8TNCnFkdl6aGjJW1YU89SFwE+/roboJBIkIvGDSJB
WABt9R+gydNkC/Soz6eFacM9p+jh1orTAgyZoHUpJfzgZK3WS9QKEJpAN6rP5zhi
VEiYkmjQme9rngaqLtBMCuKRHbYv/DudwOh8UNKQryllixQOq3E/svhBvCB1b1pw
j4ZUBuu7KIbOq+W4lpON0pc123vCPWgrXptksnGuY2kDoSc1GTBT42TWoKX7O/Ud
TRlG0leRoqOz9B5AOFgkxi3YjxKH6S2O+Y3buz8UQr1MQkuvHxZwJ5+ojerLN2lP
mAGdTm0D1rSMWMKffuT1HRuUFGdl14qigWeVn+DUxv/MBlOF/Y+X6AG76MDnJU+h
Qj4IXCWt4DSjapzBENVITAw46k6ysaLD8qJO/drLHgmzBlFhxPq0oZOLUVYPX4YA
Q5c7r2D95cSuUiryoEQTB2W9L3b++HVA7LbB1UzddicA0iDUelBtie5betesplkk
hPbvOpnkUzL4jlxnFk9l0vAM+ULYcZ+ycdB4pSUQIyVBzFP0JtvNYuKOy8wEpgvx
orMOHDkWmO5hlbHOnz3A2ItNd66jwp2Zb05jHp9sLbjeX2lWAUkqAPUF9zOPDlAr
A+mM2kMBTMyT8dUv3ai1HJKYLvP34RoJvd1thZRbao4csMl5MCNeC9AWibQWdHAc
Y8rlOdI0PQlHA7paA+MgD/8OsTvp2Yt7oxesfVgCc2/AtmrkaMlTa1rPKNCs/0sw
2kAba5swN1rHQmH1vcADVjcpg55lzpbb7LSi9pQJU2vyc7ObJdsi8UCDoDCgQgVZ
lBtVcSkfvZVTmwx5vpJxpG8hkITioe/h7++sKFr7l/HXn9VfF56AHBD4bMVKxEE9
0imU6EwISZdWipLtkJ8N+ZRLEwXyli+S/KSO5bKIa+SjNRyh3TTI7VRQBnZD2tU3
dCViPJkeu3m+/iVHXjtcNpaSxralzSbxBkyhx44HzAbR/1//G2o2z4G0Iqgoisdl
ss84nxRRsaSPq5L4L0/Bs2o6J+69UECM+4dRNPI0pwmdOpv/AROHRNf9BQ5olZyO
UKnM4nypIoYjKBkLI+k7twKn+9RUN5GmlCCKKgpM1KsQVQj2yXNwpsFreOBqbop1
ujKqxJwWDOCPdTjA/TP+fudyxE/MaiZJISpK7IG5kpQmcUtfrMtQDQDqARHNtWB6
CEHwzvDeiIXyPLxSNoGlFEnW2LBg5i5e2B2fPKHbC6P4hXfR5scgNuI82Xe6lURw
DOxNpkrcVgE5xwGyWAgyAstvNDQmVaQ1apwXqlpzvc2CllloiiqE8M0u+MYio1eh
1z6h9Szj8igYGu9JhEu2P8vY4g+lGRfRcMK65WgwglVuty+tOiNAZHzaZwN4ECSz
T/6H0PEXJNdyUpi9UWvt3xOpTugLpGyyxpSYnQu0zkWG8JrarBCPvSb1p2pjwypW
t1hpHbrPihdbrf3P2cikdIHJW/f1ucRTSf2Vdo3/WVC8dlu9JEld1MwobohW29UT
7fGPZvDS300analRCyZDM8ZqNFOFTptdm0AbzgFwrE9Ml7ANStvzkboL0Xcpldio
oevkUSO+GCUtM2Ixv+GTQbFt/aNkW2BWQnCNj3reIWS9rWDQzlnuEqatbQ2IlNJ5
dTpt0U5sVgYWliBjut7UHBw95e0L+L7qOTDAKQB9ldov5a6B1eHpCP3IkQOeeMxg
9lEeDyotA//G/C7HhsB+RCpeHhaRBIapt7yHyu7mlzibonW5rMz1AqULP+gnxNgW
9clIV6wii0jOe8I1xqWSjzGOmRLSSDWpfbrw1R66K5tFc4cDSG/ONUd3W77OXzYX
5rtaARNRthf1cbMvVdVhilt+6SaYNtCoN6GYOLOwS6XS22OvVx9hiK951xLMzajA
i1HvjLSfTRXIOYKHpR8dWBK7JV+7Mc0UQUWNpy4eYBKow5gBrgx9971DQ0VfTY39
rajF97wduUz70pDOTA6F4fHNhDi5hx+VZWOogmIFSkqqo9L0ABk84BNOOlYXyT46
kZvuZfWOuFXiLfl9n7vJDPZALdx0Q9gBqu4jyi5kuUb0jaECFtwjemqBZEugECap
EgcClKXoUTku81LUQ4YgC0SFZu2h9KsK5kegwu/U0CZHRjifWiIjZJaz8ODZSxZq
9VQ3RtKuzODdU4uU1YoXV6XVAO/Uhcoyg3LpNQcsoFRFGAXGush+FLdTlNUN+Nmx
l3YaHgi5+UShBfwnRX7gW42xljZogg1PQwWDgtD+Jl+K3+LCD4MyKS60WMz8xXps
+OJrgxjLz5X7YcrzWC5bZKoVqQTc8hgCBwd31E1JhOASTMbz3oDbiGk3KOMxQcuD
qRop/tuNPXqXGBg1lXZxMRUlwSaRv6zDztD+2s+Orzm/1PVx85E79sF1fFlkSz0r
j255Sfvc+NzWGFLERGsZg58jBTKYmUOkWVs0771LXb6gq2NTyyrgnv69OuFoWsJ3
BPzQGOBoN8KF9GLoTQg92zWWNVosffXjfF861ZZKLrrHMwTGQ4Q2uM8UYQf/iRjl
GAJABEeE99Ubb7yo7/q4wOSZhANOdiAMB9GLE6Ze9es33fkDyDblkVnqeLZJG/bw
OV5MA5MLr/UPi3ZH9Nq+I+LKSAhg7NwXvTo18ehoN+/UYd9cotdSWtO1UroKWebl
1QScKKKLcagEpQOIfIeTyEQzqRURc0XM3NY+m2XYGn4ckkHpf46t77UdTiRa0Ccm
fBDnOx0p+Ur7ghduOONQEgEiF/JGUKHi5npGz+IVwTpOQccwkEenAnYU7sMMT+Iz
R3yC4gYEgqsJDbfCcfbbTnwI0D1Nbr6SkJ+6N8bwTlDTcdiWH9RWof5LdL1UncAD
cYx0W/6MEVOfpHxY4jDeR5s9pBldirsxjUxdqP6p2vZt0c6ovprPMHFynQxlOg/4
svitSmRm+iLVet4Fwiet7MsPDeSYI26wvTGxj6/dH+s5+R6W4LShawOuzya7DOET
LI5xKFhJX8Xx6V0/rJ1Kv2jBdZINkFWf5cueqOmtnizQJh7VUjAJ7BKR1K4Ivs3P
GF+aeYOHYsUxyn8khHsEf5E5Ha3GbWEpPomjEAoBQsWLjO6md20eJ0+ndChM0wvz
KFvhaJyi1acT528Q+iRbk0aT7J+bWkrPImSxezEmSoDf4uZ+5Yyzdmmd7fM64E+w
xQrChMWp89OP71cSCD0W3LG9tl++dfBohxjV2VvyEyw4mVVj+qeOqldxUbQW2gMe
Nu2lZqQYYtTMnofEnUKMHlNpnrBcloClenbKna4dR+j8OubIH+y/R5t/qtFa+6f+
QP3FZO1qnL8fSGFVAuKKiszbPOGRl6RiBbeGjJe81vXaGx/rRiq6vcmSMGFhTtYF
75xOZHFVDaPhV6CcL1rT8av+7kCpEEG62yXIqY/kS7S2OgA/NewE5aK1/0jOy38q
lYWRsHETnuFtagrJ2pZGNt92nTNftC4Sj27lxbkkQh2wolvplJZQ9WKaH8Hnk4Lm
tcPiDAECYgIA6H5r0zP7179mo7Nmx84kjv1IaYe0A+aCe7M+twkmJbIylNEjRTvx
q5+r2aQZpmhuijNw1Ik2xc8gkBJOwRm23U4XAGKI4BEn2Jl5tpPXOlv4OXmzguE7
fjd+Jt5d39T0ATvkXxYe1ROsYD3iPO6aHftfzO3T/2m42BiH6j8YN3Y25Noz9JSp
s95wyYmK7PdTu/TwfrlS8HQp/x+TnrAhbDOmkh1w0XFIS1nrIX6bMEvJzSVxanPX
SqCa9LacOrfycKa1JV6onC+Ql3qT1jk5Mz93G+uZ10fv1qPm4w30Fn2tDpVgNoky
lGACetAIPKnqe2hD8BGuow7/RId3jTgiNfNPl1Lhi+jNEfp1jXk8053kZdbpW2O3
F/Vt8xGouuLY8P16bbZ8j1li4fMZv2/OHQpWMwguLx3e5yGrEYn5OUcRq1s3P6k/
L3J9D0NXSrDZh2KnaETd9UR0ELdt5+2JXCim004dyQmqywX3lmeAQAbO1USHfpRB
fJZO008wI5IiiWDic+1PTDMvL+4gQlopjewSmnwzawu4ZN6dW899+z18mhVuTz/G
6ty31oxA1cGrM+miuze2QprSjM6fmMkgZvThHQDtUKgXwofZnjRCxZjAYQuxds4D
qboqEtGYcEjsNePxuLoHYB7iGqQmQ0QzOUNJkyqQNX+SBNCDotLMrzel0phUdJBs
/WqCFBHzPwn8AZlNAEO/up9KYY27UdKwe1KIY8B2mRI/tcCj18JqNSZ69SHdKyz5
A7c0IpO2EbCOpDndGtz4MXyRPwDojoNmehx9TTIX/Nz6iDOweEeCXkRKxRGPd9y0
lM8v+xypwIAud/uIoIGrgv6qimyxYLBEfUjlSFZJM01QHvJ3ZqO3144mt801H3iS
eV1GBb+VqejgFsip5K8Ekvw3JJIXeqdsVUpGo5pmPoADZypWyymuNgtHKFd+xJfX
1EhOBgBuYaPxIE4p84NESgxh7BLJq6OeeI9Q9uo4vavkUZrYhsT1qIBy5lHyzBEa
be6eE8FMELLZGdliSBPqhh/PtxWXo8I/lpbG8V312sJn+zVFMns9PKQTf1IXR3YQ
YEn3G+8s4/7GQiShqDEcWp/MgESSTpHAJqCifpUAaROYT/1f/QX8hRQbD0Tr+K8s
bJw/VJLBaKXwiJmScbrAA/adGJQ5HH96580GaOSagu+t7yi3d0LpNLrIDbsgqPqB
h4Nj/L7Gb/2mtNHYxH/nIVIbMtRGa142EFiT17fJp69M0piWw8QVbUmgNn2frgJ/
STS6foVGlZ4qpe8Cku6DKDuYG+Renb1jzglS16WqBdVdI/5zJdMd/jND8R7svF8e
qb/KKF6HQabJvaf87k5suREt9Ga5gjgc5QCtXHZbJ5TKgplVg0aNnkPkHHSNR0D0
HaqJfXAK85dH+yVO04PTV/REwid4E8V7fw4T3zI9s65GsnNb4cBzYdvS0UE16r3D
f1xavFkGa5QioDA0uVxNCUtzhv/6TL0G8455ReUm3PDNHw/8sgBaHNwDCsedhm6j
EmJGGOxXn0LFHRe++zRfZS4xZPcvrNjj9M0k6mytsR40zxDfV755YNyl+0Cs9YBJ
2BDhEhL5ykoN+XSu8HjxcmUkLfw1lyZhG7EUZ7DlKwwddf6voRrttDACS7InfNk1
EDi3To/sSRDi5WHlIyhg/klqE412hKaSTTwDJDr31AcKGks+RtEFMPJ4/99VdPUW
K+szL1S4aaBrxe6XiolbFD1gDCscfzYEkr5Ybz5pHNzP385NSYb/uQrPrLOpYu6Y
PVG0H/2sPTW4zXpDjhd9h7/X/6UD+9qON//emaSWZuUdeUp5tPR9IXRJIFcf2gLw
Q7zLdFlR25GbkO4TIUhGGpmsgFpIZ+MI8elgN4DEd8tzuEV69mRiY55Af0HbIwGe
S+xRKqmOHoajrlGmESE+45oP5PFLbUvKUAXpwqOAa6VP/LM+UAko4LNNPF+VBfi8
v5tgV6of/q3W7jMbG8B9DEPcFmlGeycHBlZCmgQFivEurniaP14EAs4fzKPH1HGf
UDrldbgwn7u83h66PhM8C4e3Js4i6FLULZgd3CgVQjYPLM8LZ4EEV+txD6f9V47S
4pekv4MvSCT6gNFS0tG+KzVpOsImgB98IgdyvKMaI9I2Wc6F8Jq7kHrymkRy0NNd
1tjPKBTbfmMZ9G1YSNvfTpF2bdfT1ZctbpigkG99QpyltrQk/CtziVQ3msOyGC2z
sGF57O2NqnRaeXfRPqRB8IohjdJspEO7QTej6a84txbnxg0Q6Q7wXvOtwMfXsiVl
p67pdBA/pY4RfNNkf7GbBeLq6GG89XnneasQZ8oZep+UKL8gDeiG33FLX+bU5I7Q
LrnT4dnY5k1HKTD4dsrdcn+8SbXIX3BcMUGRtVb+dztzdIXfQ7jo3cAV7LkJulJN
Wog82ineDKPUXbGdtgeKwHYn7RS/BL+FGVcpmtx6uLEHt/xe6eHI8xzVjUygyRjk
mThfB2o0uWDrJO+pxVZlxrzuDBXheb8+7qmMZZUPrOnDkhf0CvKYSrI3dNwk78dJ
+xkdU2TAilgKRYKajOPHJbqYwMoEWwhMivm0AYI4RR8Q4exh1NaVqssx4kpMF4Bc
FdbIlrFN2KyDFbbRcajvNf+OJMvo8+xgUkfXihEv3hqD0AI+178hBSQ5z+6SXBU5
TEdaT8rcGj/2L+m8pcB7cXRncbHUsYQcgYmnccHSlDMJqxZW5/FqMlhIU0qkY2LS
y5xYZVt2cH9QlR6URSQMpiNqvxFOz0cSE9ZPcdsAFrP3bEfGFGKHrDBLCW0NJePD
wJ6FR/fh9Cy8kgYJaEPowMj768Ec0Qqd0UY/uQp+nn9Vev13XXEojmvvulS8A9WZ
opxAqMKUlarJD8+VUbbvfTGLQfPVS8HIauXqlOZVnG57nJ4RW5W0ttTt7mik0fQO
IKdQj8BoraqjObN6aOwRyYeIxULgDDcfQS7jdSeIYVDIvrBzEWZ1K1sDyYjoHRxj
C58o8jAIQXRA2GJlVH97ByjFcIKy+FNkFzr8kdhNjhmQNF3zOx9kEvcqDEJ9/3H3
wF2GdTYas2i3ZfF4RifMpoOMQ2o9a1Jr6RzPhyjkSKpqXEcuZw1lB/gRCrv2sV1Q
kf8TEEKWAtge4OmX9HB7bL1aW+/5xPnv40JnDl1iC80ZQFzt8jXos3u5difMzpSc
qQns7tTKYh0p1ZFLp38OcFyCRFJ+d3e5WCYBCS5gw6IsO9W47BBdMKAwqS1a4Im3
kVn4QOXg39PaVTi/MGgChza5946dU1L0hlWInrR3ThSyZqI/GVxLtvB56MzQIjI1
iXQoC9kQPxbdUbmyNMeiJO2UDc93v0txFTUKkTkl5N/mF3CTdVhUXeTwyFZcln8k
2WWqeWcp84RuChm/kVF66WFaDzUPiiSddL5s5PN4b/Rq3dzs7v40O6RPddRYlH58
sPoOXtIDqIT5joYG757b79PLiaOFYSCI8Ap3H/5eENotZIGxLepRLGVOIvi5CzsM
CwWBGlxYIrKQFOAu/D2JjJKRZPdn/uyQ5uH76gmhaYQdZ01NwO+NuSws5tLxjfX3
II3gauRIqQbCtrDUpFWUUiYbc4WlacaT/WCesWW/C9Opr5wkdFIFAZU0SzaSY+r7
VAXDWmF3GVLLVz0JTWqw3oICcb3OHjMon1IL46ypErDgFsCVrE3fjk7oLgq37oot
eop+2ZPcWAYN34IVbYLTongJLECkwjnM4YRTWl6+kcQp9ZHxNqtbahXHNFndCuq2
I4y15YrrHVbClU6PVfgXdZ/r6ZRKSKra6lOIZ76w/EVio04EeiXMVInLKsTOLntG
Q6YMUJvWi652yugNc/dWakWgw+WiIug8OlBoGBT8jzcOx/EQ04BwlVjzPaVmv6yT
ECuguHhiDyZujLv+zltSXYjn8rYc7NmfdgwzKM7zEgIA+SOQ8UDlFGj6vyqk12wd
noivRZ6H5HS9qo5UCJah50ttAfDZLNRxALb5T0aLJjDYA/Yo2u8Y06ZLyOFky49j
JAFsXbFUUbsZb/VbqUkZxautyEljVLwjS0uvvJ5JZSnUPcT2cPJIpmv1I0S0BdrB
LrsJVTDXnsDIG7hyryNX39GftO3alCJJollddyFssSuZQ/qnEZzE3cuQ/NdRgc9P
REWWaXfWN5ifPKjoUr2GHTEKtFYmh9xZEGvhGy9M3UcD3XUD9gvBVM+M46cF66eJ
bZlVhcyGXpo3BxUpH7XTnUQ6+GkxZBP2ARIjz/3DvZBBW3e3mjzts4zkJvj9H/m0
GjXiewOAbY7vctTbY/EZCjrJmItgOMYTg6th0mtbB+AgkxMIEaxEbQ1518wgJBde
ZHexddY07X/yDqvuO/+JxL7smr3DZYvQ++fY9P4Nk83cGVbHo7fcrwNUhL9e92gT
8kNU0/anL412krJyrLJU6ykHPKyS2sln78MaWwmZJisy/IISTpC/NrWhOnDA3bHf
uZfNQjlv/TH4C65JqSIhc1N6Q2iWBGURMYolCJTr9/WWdDqkFEZpV6F75s4oSRcU
jeMttsQVZMQjLY0mORsYocZBV75UfVBJRtf8EAzgByIvNLgEci/ebizjQqxR3Om6
McYrGKIN4YX3xXbRR9WvP/LHUAEVPIyZXFT9nLPINC38xeJ92Sorh6FjxLqT+Y4Y
guo2432yelb2JfrDmAuz+NoJKOF8rNVkRsAYDV3zHxYFCvpoSCr+lEd/M43g8XNm
NWcPnffQfZUsR6LJRx9RbPPeXitjvwPzjpn/top7T4CimRtb1+Q8qz7+yi0FiVN/
FhkLHw0749aAm9DMlDd4JUhgc0x9mexCvxSlHj1T4wafF1eon1wIH3JnLPcu0pC7
Rbi2mRN3W5fp5fw3RdYqXvVN8Ud/g2BS9ji3CyJgnzoTDgRm1Xve3AnlcIGF8TdW
b8PqJHthhwcJymBUF1ZLmoIDRSq8VFmX9eGSMGyMuwxqSlLWAtBsGajLrNM4D2H5
cEnRi9/9qMuve8V9nN8nX7iPiMAwKxTbvkKXOl88WKic9kD+9epyriJuFHVZLXPg
7fzri0imIDA1tcTveZNVpW978kCq80dlb9F7/IAPSXvR20gVViw0fnYL9DAuAYYy
z+UfZtlQZZzc216K6M7VMWiijs33Uosbm9gBUwmHElxiCoSyneAzfFKiTXn1jTZP
TRhPyFZdfZZJbPdmcCCOTmwroOhd3bS73PGdpWqH5AI+UrZ9WFJbbfrRV3UcX0kA
s92qpU9/FCO9J8JH5+yMMdHIjFLiGKagYYKPtj6J41onmLnSfGeFMJlF97sHKIRK
iQh+31mwShUDEBNbjs8Kos6A98TKoPvfon+VxTfnBogWu2TF4tDobUzfYfTxn/Bq
QNzfgYkqjq/7p3hXy/pVOylAavcoX7PL1AaGmyImUEVQjIB05n2gnXXgRKevuyTi
szeSQCJagPEqkhYBuHfrHA7KFdacYeBgLkheHGw4l0AIwfVWPq8+6Dt/V/DL87Bm
HLyYNToHW/ZGOx6BJ7EHUM8jmRWMatB/SqnenJcst11emEduo1aHGRoFxqElLKhq
juFgwfaLOWHzaJay7MXDT2Idu1FdsSvfOroSxOOAPYLANO6/1lGcoJNuc9alXsHC
o8oOwiFSnvdD1XrGZR/Y169Rz6TDAiOGUHLa5r28S8DJDystaxVr24ELh55kziHn
GZ0BFlthBVEq+ctxb1MWG65HCpgSdMi0lk5Vk9Pr8CyUN9AZYuqbfMBTwufmY/4C
RC0PYlFuHddUkTWDMbLnKR9TQII1RADQisDmnns0zjGPbtrgb9LlWUrgWhXlKQET
HFB6rEGvtckhxwe1tIgSEaXb+xBJ7SZMjmT/dhToolv3fyd7MHlETj4LqZAyTDqs
vxNcTWw+ZtjxH1vg1afSJAytyfzkNtcFE2v47jMI37l/Ub10EJv66r2DpNjYjFa6
OsazqH10ddwL9Wj+E667GpWxgJak0HH+nnZdxHwVhIIP13S/svPeS8Jd5Hw9KPtE
nDw5ZD1KSaOzSxdRGsyHEm2wBiHVGVqXunJPfraqUOhPgHzf0UCVQCHsMtKeCL8C
cB4EMUeDEqO1GenE6ebzeEnaUtBfURCnOzCI0SE7jgYtgBVK+asA1Cc4XvhBxPz4
BbLGoHh0omcm/REEMld8ih5mVeKWShRZMr9DXa8Ld2xSSTUDQQ418Ui2QLYNclSa
WqEO41vkIxFCQ+mszmzc8cfKGLJuExGiBN/zRsr58dRauaButCrk+tS4lRZ8Jh3E
/PniAb3R82GqEJyEKKmDX3qx+SKdpCSZlV4EuLuzHgPEJ2g87pQz7WSxJ7gJmtQT
f5PlUcQG4BFj/9LG7ShD2SPMPcf2RYeZ6y5RNWPd6r+O7j5+t+uW3IukZ3XKGvo/
qpKOfymV5Me62JuftqwMYHv/ZRZUPsdmhkAHY3+W4omOok632C3lqsjKKuxeF+qB
HXhmw1WqgZR8jluEErimdVTKUx++MTvNCVXf8IqRWyjJlxqrSPIi0ebIv5OXzQVF
EPgqdAuf44wtkvQ4cXHfranek681zQR64HBbxZU9sq0GrPYPfh5DjHZbuX/+ctnK
wUQi1c6daS0Udkh7EkMEeZTuYfOqi4gUpOe/xmT5FRol2pSgWCmlIybVWQKlmU3x
Oa8uUEfNHp6gS9QsJe+vijH51x0OiV3GxzuzdmIVtV7dJDywZPS8WV+5O92UvK/+
ERXJBBjU3niBdIrD10e4pw/soetrEHO4RMWTpwRLB5gEIEvzzbPD6OzIJgWYA+XL
3OJAZOwOgiHS1AFJIpTEYaOD+mhAiRoeTmHDfnkWkFRzVhEq4Utvymogyssk0wfw
93l+HJqLDoKeNntIzHf8gd86ta4X04FWXfGsnoAgFZrSuVxPX+lOsNaV/FCr6CQh
y1ngdOc99ylM1h1AgY04l4KUvMKw3Al8hqqMniMDbt7t4GfG91Gr+5Yp/++8Yt+p
hjY3UKQucG8XIMS7PVNL6c6xfTT0S0itGTD6Va2JgCh86bxNjvb9O0h/UHO5aWg5
FJZ6MFWPp6cAMR0APi1GBR74fmty6QjwZ2UYD9rUhffADQZ8bdInjHp+famEVNjR
6uCO6t6ppVxPgJsQ37Crq0SmXOovHW07ymuQWNEiGR8jp2d7PqVF+HMCPgnAZ4bK
lXcfU+24k/Q/Zl9hM+w1hj674/9sifwa/g7kuvHRkoKOAC1ZrrMq6ggAc8wZrPiv
7yAu9PUzflV2BZSA9Gi7RxEFjqy+Aaf3jIwjqAmd7C6uQDj0Kl56zNeHiv1evumU
Lr8li3hhKDQD/Yy0pt6GDn/j3y/W2U+SOb7PBsW1hkaKEfwUYaBdP/XBTAX9OwkG
wSKWTG0yo+82OaqQwI2gkVfFXNowxCZ3cD95lkES1SdIhakTfKkMLUCTU+J5ApJH
4xP8rPlVHPvMkix5PKDoKDZMU100NnqWJbYjB5KzBi/sFunlvZvj4RGD7h7qQsGO
uJDBXYjhMlAEvBzWn/Owh1SxCSyebIA4rEgFOFzxqMpK1QmTsbmMiZcRYvs66OlJ
tde7T0JOUlwXg+yl1riaLTtX/td14x4/169mE9UIjAOVfimJ/RYrwKKobToWrp89
lKo16ILScoUk2CcgNZ3C59/zeJn23nejui8Tt6A06Rno74XRB1xtTUebTUGNMVtl
gYMmYzxnaJtSnyFx99b6dXutrA+yZALAJaHn/prPNknvMrBpQrZXiiVTIZQEYSi7
4Oabl7Ei5SltPvjyv9a5HEh8fJKIwzrf2QlaGKAcHFzvt1VsrBXdmYMKoIahg7WK
GJb9aiKG4DyzGEAm9cNJZpmzLEnL8j8wDw8WglTkJavav1fjecu7Cw8cpHDBT8/X
kkizo83SAM083y7u316j2rbPCoMp5k+lD6qv45N8NHR6kXGARA7h4SYsEOb7X0/m
N+DRUASMfJryc1EdvyExoZLHb1t9+nDpDn4QjRC4ZGXypOoMQy/Iaxtu+BOXVedZ
LX2cfBm/HSSaEXMiXzLuXtqf3PlMihNOT4xrGqdga0ZyVVsMO/9cXjcz5Nq6LPS6
IPvxnVvd0I9djoX+iObWZrwdGBQyhmJ9ddVQNJi5WKMKF8IWO2klNkv2ARsBNJHf
j1kHdsPkFP7X9h9P5e8y6sSeWLF78hg4UrjL1BxxHexXcUx6oICYkCUr2/P1qpR1
khUeVaePpZUHzP0iVT2JitdWKW8EZlMiR/049QhI5m1emVsp/I8mkQ9cfNWAnOPJ
4mvnN/adQwn8TtbO/qUZdzpdJP7bv6r1Z/tFtiri0Fp7FN31wmfc3skI4sWXC60Q
N0NbwAcmPaQHrXjD+8NaX7YQr2Xiteo4wbbRYqVrEenq8basb+xWEj665nTVG7Fv
OS/uTCPA1i6MIeFthYDCKIn7BYhTup9r85da3bUm9gLDrm7EqceIzOYOL1VE4F0D
4MXB7uQ0HRo5caF+SFfVcEIeZXA/zuWxp6CayT07p+lF/tfybJJOdhytKHjv7iaT
HPgLYV9F0GxNnGmJMFIAhoGIOQdDCtRLlBEEHGpj6LD6RuRzMPL/Snk61nq9JUeD
4axKEi6lwneUWrhdsEGPszIuwXex9Ek4kb+n7GfMSwq85EF8l7czUvII4MH3eBZf
MpSZF3O7ys1gdLMxeT4vykzZLyyWEl7tx7C12B5fbrTALrGSaPqTuSFinQHqNIlk
vyNCBgFTO04Xb5myEEVHra//hnsGC5EteUk/VUmNtvPFFsxr0W1tMyIIOubm3m4b
AuttfQXpJD1vTU4ZqvyRiwzrowtMn7zZm/yVHzl/hgQnx+3d2wF09XmZZrLL/El5
bQTqHAEDUkWiAE4qPDOsqdJKHLiUJTxld2Zzm10HNEnOZUD3kZpk1YFyTd0l30uX
tfQrLTj0fGs3z15/X9pRAhIFgHBNpeVKy0SVDpP50nEKCwhIsd09ZGq70fef6GDa
m2OEVmhcF0ZLatCQnZJhD1zlyo3TLw5ApzbZIFbuEp8T/mbOfFCEKsdFvJHhWxt9
oFouwxGNzDtZwp5U/ayes/zgDV4P8Jk10eurIuEVULKHXd+rdvtd5Y5uFXIGVjFt
nfp1UuhlnT6on5KjYZ6XYNC1Z7X8fID2xo5h+e9Pn7kdmhQaPUwAUYj1B8ecMwuP
7LcKv6LmKYfGRJK+nck2hC1v0U/atdg+/7Sbt7OZ7H9nLfuMoxIQ+enM8JDB5HY3
Uv4RKdmYxAsH9YoWEkSCJgwhJ65elN2PtBwxV3pMamPwHPUHPolEAkKZ322AWp6y
e/AC0PhgO17uX/1tQ+KbvyMFasG+Q3eyMyL9znj2G++Jk8iIVw5o5h9KKrsugJpX
gNmR1du4HUlhl1V72FGvmr3MObsxKjkkv+He1gSbjKwf3JeGPwDDovJJfOjpIiTU
uxK7PM2bUFfKlOxmETtbMqEyej8XnyFpexaGOITpGmqypUoeUO35oUFr/l/7L4FA
CbtMYjhQz2VHE8TAq14W9TpVcjqL6ddlMHKeXHgaQGoNFzcSMLGten9HMQefFpvm
m4XdnuhLZDAe7ZoJZYL1ILn5j5CMnGLosvTtHhJA8ZOb/R92vxO3KngHDDqb+bTH
oMBReTiYwESql8M/tHN0ZdXQjlPSVT1m1X70SJBpHOJZwEiQoL0Wj/NWfThtcHW9
ewhF7MM48CZWKgWarqIwlOI0non8kZH9K3dH6aCRUxCTBIeHzoC7cf+Cg/Iu+rCE
LBQiNr9PQjnyW0FIdvfXviTqTdNlYgzcTL1IowJFJ5Dc3YVVx9OTmoIAdPTnqMQU
IuUExgSqjPENa0SEmzOou039DMhuNZmGdXGQhcYxrkc+Rd8Iu5vL0yzF91QDER6u
/zfP7bXnMtEBSWbbLireEQXlNsrk8aFaG07iBJ78wzG1ztmx1cIgKULfhgOTDXFh
RbvK3mv/q3CeZfcj1k2Vol240w+hsyAlzitTLEfvmCLSGsi4NIID8C5DwpOiewFt
x0ETXe8uxVz2+f7PWwsNYmD/9MzBXGgIvWraI3x0mmpbqtZnWm0nkguw+oebzKzh
yjREC5n6ALpiGoASbr3TDVLz4ES8RUyuZyFksJ0r/OcRgq7SSK5mDm9zWgANU/Xf
EUkjLFxB8jrXaVNWpip6fmcg+jYWPglo4M7mFnOlHr5P76VLWTIUIbktmepNj/oV
jfYQfj6I0aF+kADUyjDtWR8HvfExAe84pY7PJb1tykZ9Lau8P2phmsxe6UBJkX9N
G59VqmIF1nUlZRm/KbSDV8Yhkw4SIC4cH3mWBSa93IPPKGA6AaO2llr7Z1Mg4ILF
oxF0+l6qDU6VEtzPdVH55feQU3dnQGgncTJ6Sc4gJzuWHneJ45mg8NTAvUZec5aO
dtO1mtMIXvsO1wuc6kQBs3MSq3CbhDQ9miRkt18HLAjuvFinSJ60trUTPsmnfAWP
RAsQ9GW+tgR8qPcZx8nyO+nda+KF1dUPe3cuGPMzQLnutUCXGpfW0tGFlsu02Vbo
KAJuYFhnhiNAF3+fs/A7ejTVdQ4roEbrcdMYDhM8PaQOIKjrsnSbRbtvmxqykq5J
H5dZmdeyxP+Mlfw87uS4drL3bhYc2foXG1B8XHREVZSLKDnxgU000S6hJA1DErkG
J35LA3B+kMyqmtG+wP1b7CNZ3HZEwmvk/5ow6y7p5T0lfi8D43sBHzjJ9LNx61wF
/X4F4NLNOyFOUjb62qs9n0KxQYm9QUJjNk2WT0ojQRlZGzYoqBLK/qJGi+bt2Y4g
YaiBk5erIqzxfPu8H3f/5WN8m5iA92hhIdu386NElS9fKq25FW8YU7RUjk8/DwQt
acVGwbZXEmtNUE6ZgzqIzp0ZNeCIyWRg9NnlXxysvt4vp7RGWa7IjkrFcVmyjk5X
dzL/11ib8k8f3HNfLai70Z2i+XAjKaxNfAE35Ar921sgSvXPMqBG5cN0znwMzGQr
Vy6vZEAjvINwsFOkbjcVCWrVYYBLhSY1Xl7ys28m4bPUJkJZ7RMJYkL4jKO2bk52
im5s76JFheuefl+qnxTYvy19bLpfxpmN/48xCL/eTjuzykL8vet5E2svQ2WW3gL1
8N5O9iyAoBEKeyzyNOWU5+PUBg8+BcL33VOv4FVAEbLmiUp//9p2LOnLynj8GCNW
xYrPyZE1hsfH8xoBBczXX2X/Xvt0Ry7LuWyu93cUYTHy99QI+rnl85VIqdZIi7Rd
B7DHLUxxJ8kL7ASY6b7lwvF6i2zdBD/2IWw4K2EluIEPhRPIrpPDesJeH8ko4/tj
XUUKijVKotr9Ovhm/u6jF+YmTZiOcODq7u+90F/N68Ab5I9R97aqKrqrzDMWNolf
uho0Tkca+3s0DkzigeyCotmH5kXLvB5bwosIwOMy6auqmsi4JoXmTsVb9zANbF+7
pTmOvNIQH+GPTHenVlq0LvebiC1W9uBj5zEYoGhJTK6sm9/W9tyM5TBGaJZr8i7w
e8dQvDaupirE6u0JS5W3WL2uYgHrlUXDINVpEw750x2Ggcl10yQ47Wqq4MvlBPKx
KBT67qYg6C0w8jGaKSL87QKFShn5rqMabOPaBU/z2isvjn/clm7iWC4hZzfwjeuJ
bwP6//EJj+Rb2RXO91MSW8GS+wG3aSK2PJSCaQd5bIF8yP6m9wk2JyusV28gxYlS
oqw3ohe62ZF30QIB9IkAme5+4u/fU4Fzls5knqo74bAGKi60fzxgupI/Ju5yp5xy
LSdsqNy0TTn/DdIySxsi534wWWMCoUnY1OunJBVrdHOeYDe0mVwcEYDnSaBii/yg
WhTWMdj6pQ3V8GZHinAlArtXp6HRN8zGox7ih/lK2pmnGwD1MI68HmIY7Wx0WSt+
LNQHZNdeGh3fpy5ZdZURK9jRTiZ3PigI95/jb9gZBhDR4xgVWl0iqO/8Sw/WE5lz
8AgX56stnogeGBC8qy4Pud2MxUwMFtcT8+aUx4Bf0RvobxYCQEYG4oiepzlJVZxw
WMQiiDP3TMAWDbB491GvHX0E6tYm3Emq6RGqj14+u6CZkyOk991F7XZkuuIRLI7C
lp0sae5vbrvXKiHy791wyvFf6C5JGItuaktKveaFKCbqxKfdEbJxhf4S+yGlY7LR
Wv649SzBQ5zrf+A1qE47/b5lTxaIOt6qGcSwJuntYqSGIpi/v0lHFTbzaV/ZRswT
JK1Fa1tOY7KGM98gVqhSMf9/LdZKBVEZE9vO2l37+VgurJxOm5qUXTs5Qp3WvSnK
fnMLnJZGY166Sc0QKpXyFqX5/z61jg9IxoC2r8PH90x95v/pey5/6w6ojO31XJbs
Cuc5QncLuM7RRa+sPqE+Ica42v3wDsw3Tmcel86AgnLzNF89+J4H9nUHSYcMT8ba
/hQdM8OieHD8Z7it1roqfBKF3HTVQDZu5sqX2p6DT0yGkOj1HJrSdQ45lvmgmJKT
Kb74P9lbRkFyfcOGjSmYIebO811mUKCpmDs6ya325YsPkcujOCrMQqRT250gkl14
OqJe5jAWfmjXHpUl9GMu4Md85O8Ytq8CjTawGwwZoG4HYX78sL795qXkOT+AXr3T
ZPSTLXvHbFB9PfMeUdiLZWqCbiRFXT4G5OVv6hrMoELyoj4ohl5xV2zqBzK3otPE
IEYagT7eKCCwFWmPa2RiYKYZJm/6foRScmVOk77ovmaEizgiNXgRTux6LVOhoYvZ
0+7foJDGIA/8Krdabmmk8WEJC95J/TbHW7ylr6Umrrzuwt9HPbQedkl/fU3MHie6
ByL3ZAHwnvtFU87XGBhIEn7k8MJgtYQjtRCrAg2tHRGsn37rwpSK5zbTtoKAUP/r
biyMeRxFng/y0hifeKKLfLLb2Gx0NLIcsWw7DOavnqnrBymiLJi6OOZP7r3UgLqB
UKX7ynYJl2qsAObjIOB13wg4cx5nFjUxRtuNDnYg3DEzx/aZSPdahNwjaeSrCI8P
d6x9XJ8b/u6IefkmZixxVnP3Ux3SIEkwwSYm/lly5dBiMDCmEy9NNhoTBi3ZJZ70
8o/5mV9P+3BTGHI0UfZ9VNXuqTlqUEAldkOm62mYFMuZv737c7/dUN/aCKMcIxlK
Rf8M71dIePQUqHjJEsuCQTY6oijIggouR9qbw8dCUThEx9pgiBxfDk8qu/YAcBte
rIuPadskyU8yF4LbcbHfL5LRYcRFFjYQPFamH/6rd3pbySNrgilo6xQHFHlwoAYI
hWjov593iGMm5YSST1rpj3628xV9OS7QBMjDDatnsEtUsa98lgezilLx0ZiPPngA
RuXYbOMJBlUjZm8OBg4tfnY/35G4FI/6+KIpBrpkmK/76KaF5teaBq+qApBviYVS
7n8E5t/LhoApqWDnxz5U7fuCTECOeUt49T5DzgBlGysdSSlcS77ruyuO8mKx0Uqi
2zJQbRdwywMrF9bksiVTJqodF8Ags93GWnuIuzipQrVX2iRukWae5Ck9PuNZ2LIx
RXnDqNVcd1+7U48eaVqFe4m5XKDv8XgZ7GKF5ld8ND182dC8a1A2i73Polw9TA9b
8AKIrisgN8+b954jeidpLscuXYP+kJoaICMrTcX2+4b3u+aOyKXnAkiLLOFvqTZM
UmfthFLPCcTWQ8c1ElQKEQSnZTQOV3j9kK1fb4/kj4CZ5Q/QYLXG/g3CL0+cLA1i
mN3uoJbQkRf6sJ7B7vU8G06vj5E4gqmbBF4NvEd7GomUkGtTcyZCDJE9w85JZvNq
jNmqE5ElX++Bfpe4DyfrBGf4ZEmAcAmVlyDF9xTs1mVssVNtTCTnh9tGvdEsujN7
DO8hiJMTVzOiSALBKsJKRIBF7ZsW+bvVLoGGT0Xx/0IygLZ1UxnW05LF1Sp9A9mj
KS4m/ahlMvM/dD/ocOXCV/C//s/nvK/iCCDEJYuW+gX6dbt+QxBBwXzpPUB8ys5p
W4kX2s+mq0a+0YkDoixyjqY499mA/l2azjiHAGr0EAAm7xozUIfKCdLjw+shSIhx
RVDxZP0oPfsD6MUtvFfdGsw2XBsxmUszUcLzgBdZKadWeEkqGBZc21iLii/zMFOJ
HArM5T0S/NOLCuN+3wasWbaWD+hiCtB7n00yIbLc1GeXqJMIGB2qQ2h5UieJJeY4
mT0zdpPnbZolFdxfxRPxZwocXW7KYXvTUeh96gKQv4Pnut9TbS8NFMXUs9ssQ+NR
8ve1gH/g9qLStBAuueWb+28L/dITpdQazBy+98KhWiOoGrkObSo7i1dybZA6I9f1
rTjSlLHu4VP2zLiUjfZDcdyPG/LWIJ18XNVAqywyk5rkcL3J/8bnyKhshvkJmR64
AEDb2/O1laWzNuR1a8C5iR9xx53g/AWzbjgAhaRey6bk9muwQMy/6TY4e9P9nsmQ
e2otDfwigbctFDMKfMd/iuozExNEN/yvCalbqzuX4f9S8tv2HoA3PqN+MXsnFVBw
n6OcrQW+frboNVemB1jAFLf5CMR7zvJOmUnRP+hPKK3Sf2ktd+BzjjEaAqqf6BZ+
g2Db/YCeLtcccwAV2KHRBqeZpIRfEl78aBqSwb9jv601ctTzc2qDRqqLoARxIMrj
r9SWmjkvN0RNQFJxoSstI1bBXrqxrJQq9FOLkbyc1/AWEynjo+ACidSOaDYtqA7q
E+Op1tJ6Q5e0J+lQeVGM8FHlc7BBIx7U1BJB2ktJZTjnUxx7I1dD9ZNf/d9wFe8m
1Qi73/V41vtAC7bUYkgN8oEy2RFr/bwAwA7uDbn+1JiQIF2WTbSd10oBgfqzRgYc
FzgRUnYqZovrpHvIU+G9G2x9LXE/Pnn4Hl5FeTZjarAeoqp8u/LS5eE/79KQDMoa
wkzduV9xw6QVMWxibYklvmLOmv4XahZXReGqF8oyQZpm/OFIXBzox7a/a2gLpBI2
xg5Wm74g+IVMrzM9zhjVKwvxcrHg9yf4nRxqdaeWXFmpbVdLDST0+P/bhbLQXeW6
mKwJaiYFqL4EYIps9E1c9ta4w8jD02d2ZnzyxnMAMfyZj0TFIfOKPUzabTDGWp44
nAHq7C7nSSoIYMfa8BmDEkQjynTHFLRw/eGMoaCA5J/iUVoExvEOX0t34vlpJVcG
GSc6ctfEB1CtSDqk0GzWzVH7YtyHY+ljN52vWl8r8LICa7syL8P2T0JaK4pCvu3B
I+O2vcBRw75aGE/O3O2o10CN13czGtXCt9eGwIni/tOWEW9UIQbGv2MNpikBxreP
TnCbKvpfIRfuKUNMYYSLHtX3+mHySEhyWIu7SMCJ7lhpG1KU+ohp9qon0CpWEetL
LSPPa2V2riNN1zgH9xOSTNs52yfQE6kj+KuVlDJS3gR9Y8sDjXPhb5x9Tt/UeuCg
gowEqqWluNP27ys+EsVPFiKw3M06FnoGw5JR8UuinmwPjOgTGc+7w59KcbWCCp8S
/++YqjZBTujC07+HdLj8C8Kc595ZF70LbTI0q0L76Lu7kV+e2kba7eO+9sCFNmLp
ElamNs41Qdemk65p2fAAO45LiqSEh0JxPzWQ9x7u89s8ZmVfmk20jfd4pOlGwakv
OwL9ipt+Ya0UGuVgVz4PJ1w6+Sc1F3k5YYDGfWHIpvJxRr+VJsFaMgfnGGsmPau1
Kw+xbehHCA+W5CoRKnIDPnGkbxJex6gTOnj649opTsBeAm7EXtAT2qKqma5M8r/H
ci5pZQYlxHeWepg8qUIyqdbsuk81Gr9jbLD5GVsfcK7NrFAx8FB+TYn57gwhwNKC
LTKeJZBcgHtOhHs4GEj8EmyD3qrAS4TCNAa4kosh4y21aOj3q9R9vksjHsdhES/b
xs+FkoHH9BAvFS2RguJla6hay5tItP643vwBHFJeVL1o0ZvdZcj9LFoVAHh8kmch
eXTCi84LIRWIFbiVw8fyidnR1yNqCD/cKMSLDUNTeVADiaPckEc5XJwC5SrIk1MQ
UCAXK34FSHE7XKPr6223a7xyI2L/g75XwFwM4boAcxGM3AYg9k5NagBR+9VeFkUE
WRomv7k1Rlr3mI436o4747RdBqW8dMYvleiqUNv8I7TJ2HqYh36Wdr6uhlRWnppj
fVw8tAXRDIgaU3bclc+G1KY768ae8iZ0ftrfSdtmn342brHlwWjYZ4ZZKhq7aHJe
RdztOyisulko4eTAmF9iCrYlpSkCph9D/sr6uPdRTfm9DtSUICKY+SnXTflhrIfF
RsN6M+9hhDTagPpzGRBy0gSIO6z/YyKScw1n8j85kAEl7+5VkIkNUlR/1G8XQXyw
zzpo5HBXN2QZC4xXF8JWh+//ximXIX1YZoWtrG3yhCdKa2paTqD6aURlp74RgkjO
xK2zqbX/c8PBXYJee/BcLhBCfNtbmaNwqfoi+jqzF/mtbBqfuMAc7zYp9zp40cCR
UtoxZZ0onoZuQDr0DuDLapQ2X2Q5xpEsBSRwYa4dr6cSYJ1TSu1Pm+5YAt4qF7AB
DsVNMn1cMvMz7BNrADkGPCBg67bYQKAzLsElF9BMhFvvz5DcEICtL0ZhzOrKjx7d
/6sWVcNj5P3twP4FLGBh0lRqYk+GvYkyN4D0QsTHmtRKKyKegmElrbmjVasoWJg8
IjpqtVkUwn2im0ybx7paZHY/MtwrssxdUJIX0ULdf3ijip7+WiQFThH1LcwcRgBJ
/Mv2pTcUsg6sV6Qg4ZNkCDBG1IxR9bohlmhrAlzlNAKNauh2Un49ZlhkB6pRBizB
ajaknHviQGe3z8WP8+uIqtKuXxgLD+ZXoTFvN65W3/c1qhlFd0/72O4TtLFWDfTN
8m6EaPcByof0FSwXS9QyZY2Ta3WdK/NuRQE2LIkGLHcHT2hSINOPyD3ZuFLSYxps
1L4C9tGygjbgQaYcn3RNqvm7a4SpsgYu5t4BqyOKD7l6FEgMiJVqSZHQFePdOolt
0JdVZBxI6CaorYfp1q4CzX/Kt/XhowBQY7Y0Jj+p0NXrJHH+tjNAEegVAqTIlFQN
hYpmDlbEi9Zo4VHxdeO956vXiv8eb3AaHA1/RSBgPUYz71CApLXEtzOYxJ6580h8
Poq/52bJjGkrC7+MLrgHCdEIQbP+F7kNTBc5eTDk4DV0gIcPhJxDYmVKYyFE4nWj
oxu7Vy/gYnM0SoqsZYE6wtykwQ6scIKM8yA/FWfwW610BULZcj/0BS4Ipl2wIBbb
kW17OMx+UTkAtj5NvD6kH2K20vvebVnL/b4Q3fd2FNUUkPU5SNszjcio9ed2P/JB
Bs/eEDrXL7dQCrudEqu9wFgq/5safGY4S2IuSnQO2fn52j0ODn+Icnj9KUXYSGaQ
BHcWytphWHo4OfVEaCDcYVmOmh41b7WOSEfN1Mje3r7nUNMQyiTIjqxRSMRZ1Rzs
o++6XELxst8I0/bnyThIc55OtfW9ntqoLRN9MVVmEwq/vtCcO97AuKY6KkDJ9ZTI
EUkl90hCAitOUpBjM/rDBmTsdAP5UoRTE8ih0q8ctP4Cwrx5aU+Is9qTIy9hJDqq
mSG0lYrI9tXqGqBTkAIpP/8OwPlqjczcw4NIF8NpZnkKQdRiz7itJsfjOkMWsB/q
if0hAnBT+BgmUNGMR48EI5dkdef4J4njvDsJBF65P0TuwcZvFf84PSJ3VujW6rzZ
huLWH2Ogpi9OyR9aUhAb5jrnVuSXV3QY38Up2275Tdpwd3Dz8CM9/8jMm9NyEywr
93FeX12BXSHQgG9hOhKlGW39xYpja8tFGf1PLITnSYjW9pysVgBlYeuQfYtgYIb2
G1oexNELEUAFx+Limn+Nf1LgCmii2Md8yts7f4BpHhWwI2Yl3g/xaBdIP6Dd/jOy
zqlWPBvKtkCakzoQaI5bBnbV39xQkOxm8SJWNzVaaHPXwyOhK1rZBfqoQu1Of6yq
lV+86GZVRDK4rw0TaK/z1CMk0E3pWxokpCnxyl4aYj7S5yAYIebE/CmUvWmwtxTd
ckaPp1gaEZ3Uy0hqRQyWhOcwkReRleJFjMitEtTFSTaIMQSS32LcWJWVsnp35+k2
5sqJQanJo/NbROnPAGyi+HZaxf/NikAVbfZcLq+5AMs8bzkkKRRaZDWzVRwoJafs
nV7+OBs8CAdEhLI1CTmTGHsy2EnvwvP7C2VWm16qgE/1xyLy/FD8txazgZTMQ2mu
2eeCxGSr6HylEDMJ04zlMeTbdRig77GYbsQwgHOLCwEX6sGT9SCYK7mFC1QQQPct
W6n3NuqBMN0dOylKOcQz+9d5mxaXSKBGcl3/c/wV6Fa8Nxibu/vUso8ULYC4wjKY
OtYNqIL+f/g08pM/ZYoWtHCnuXQXrLMw927MgSD7NAqrn5hpv5BzmjC6b272R/lk
Xz6ZjMpyU90m2i2F9TqBvYlVclmaGX8+Hqi1aEh6Bm19DM2Nm06CN+wlP2XVrahe
wvtsDGZX+lWIfhe4MW8S0seBmBW8weBrcZoXmAHYSMweFB93Fhr02n8Gl9sr+Tt5
/mHFhAf1r88qu8as1+0Ve3tnwuG8U+D/7N630EQBvvLWU96PDxs0VeAHt8X0WL+I
sJPT5Bs+5cyDo4TDXbePgd7ywkPnTmPJzKGESVl2LMHuBWzJ/49hRxH7HG/cbFZY
LitOr0Do3rsHQX6x18TRFo6ek6sMCoo0KlkljQpJRL60L2XDzrVz8f5Gi1gO6zmJ
pCOiemhemokD9uji+OsMV5+zQFvhuCE1+4SI+7ilNF1g4dCFQ+2145F43uY90u13
iAFUYBSdDPi2YC8fU92xPGrJLeVruoBgcxvwnh8c2t4jCfy2Fe5a/RY/JHJx+iKc
PeYcNuHGr+n2PgG4gw49eKpD5GgDc4zg8/Vj3gvGMH1fzV3z0bYanjLd3Pj6Z0bw
0rQ9xTyRLziZgjU9ltBEUywlMyNouSHL6tMxcYP4jxBDfE2T/HiEy9vOS4kZi0s1
ew+dO/cfubgbpSiXV9Z5kghkeAmGC6JwRucv8yzAJObbiErop1mW2LeOruiAq/Jy
INenLdvth969k/Zok98cq1w7ThSfhqm3jv/qPHlMBiQUS43l6rabLRNgVazMv3OB
RbF43DkoB5B8leNL/V2mly0SJzmyIrruXeuYybKsMvJI91V3v7Mf7YsWe8cTjLuE
h+C+6VKtvn0+mRmHbMqx/nMQqNuh2aWBz5KVmbT6EHA1xjGSqi6qw1Ax67SP5cFQ
/Ng2iRLEY1sOQ4FdRXMZZnJfmbEVnPyWYnsWBvGn/XLN30fepXer6ipOrDFHmXwk
fr5ElT9jVb7bsXYicc9qyN0FTaDJkLxBlHcXsdY6+lpLdgNIoNsyVqOWoejMv6sY
1z035L80w1YeCPqTnHIBuoWYFAsRnRIJLfh1kabj4emDaUOru0cIa17mOywrpK7V
LOU8IaP1CC7yyNzyosqGFSKuTk+j8iHz/t90jsbbDEuVVW3GK4zK7G26vpH+On0J
DevGKjDWvZtTmUmVhIV8KogJkcQZMwdINStUZucLhyxnAPxaXp8FlE+xsnvJu+1+
GZZcL05Xf4Hp0j9c4s32e7yUxOIAIrMr+bDvT0kTIQxueK7j/jAOGLYgtbkrQ+pC
c3X6+kc5oVuCb2knrdE/qRodsyFpRlpd+6ngJO/5OWF663bGXKBjoz6xBQQf9lpL
JwrpbWIGclu0DumdmcnQaKocWHyCAouhaHi7uMaNzcVwcNwWdGhuqQanxF9e3hoQ
1/zmtRPbA2oSaiESxhxymQDRjGb4zHfTJnYc4rKiplLBTjHPCeHbQ62Qka+La14v
AqyN0jv5GXk2Zxa1eR+Y6GPwHOLqyLuSZ2bEGz/D0CjCo2IA6Vb/ppMm1jVay8cj
dF1/ppt3G03ZtU62cNbwBWa70r/4Ci0DtBiJ40/3UStIZrGY+oQMScfRpSAV1efk
PfDq/cmwmB4F+3VXhL7olnel3c1/qVn5UFzMI6HXxxc+w+LHL4ybW4ay/iVeCEvB
SAOLG9FXhYjwpna3eenYuDVWpzygqNRNN4vUFyQIhHCftY0RwvcVm2PGE2FS5/oo
VQhlkXSTKhhbBZg94sN916fjnWqhH9kBNhqGO90gVAtBzdioMfq12fwLSnG3ehNY
mUQ2E1fZa9OJP14kFkF9eJto63fe7nxQNyFoY+5W5SDr4cIqpEqY8rTt1t8eEHU8
SFqr95FU8gJmCluM3a//jir0e7aKn2T7rCE0WeYTLZFTCLELN4rdHF1dFIY0Zqnd
+xPWH2hIu8tIwoBiElUtja8TLKTUgr7H3NCNYXIVZzSEELIjXBmfp5FizylYf0c+
16CII5I5aSDHHG6MEM3ZUFSiqQnzfurFjCZnEOCkVg/axpUdW/ZvzYrKrQxIKAzF
JULhZbcWLceHqHuMeAXUEKj6lZRv+NHKqUBanx7TKJnJaGZWxBJ7lIF7sIHAFEYl
9gJ4sBC8fpkhJUQw7c+ygCa7IgQCq+e6ebzGXWXJg6/klPum6MhpDJph14vsoWfs
NxXFAstt5nIBc6oLyUrrNbxPI6Rjyt/CuktezkvX2bRm6qnnwxhEtLwvfDsAlI+t
jAtpva5ClURg+jMO2O2c80yGeOl8ULRtZIPVjCdddj4HRIQjsVqa0X8udmvBTfhI
baak0glDCwwnWKYb3W/9KUgmndNmZ6kRZKzjOB+CyyCSJDa4T/tThd8trMf7MYdA
nxu/mY7lvPmUTe2YxCO37TNFPnlM7Uc0F4LogItgNnhOF+HasotYWy9D7FTbUdIq
KkaVLuK/5a3RxhMKW/r9Rj+LJJRnQEi6wvvreJd3aE6tsiOwNvJdmV/ESNE6WAwa
aOXm8zilvi5Nxa+tdwf8yqJTmWBXAzvfJWnv7rPwW+ZszB2F2EXibMET6T7L7xGc
7MCa5bKXS0idUwIgUu80eLG3VDgRVx1qFE0Nh7zTmS/wKs/LFilDCjFp0b/ohCfq
g/9u7P/KipAB/CpnbRqhXlyINMR7XoyusLbQnTLdzAm9K/PlEQ02i+ZulS0wakDr
CRYDBGCGl3mE89yFFmTsJAnQMZep3Yt1ita+cP5niaASAH13YGn4kCZcp8qdk3og
65zc8AKNuPzrit0FD0xtNW+DB6qEVeVx6XOfxO3/ToeZbZLfoy443mg6QOUu7dPf
RfQD8eyfddvNXEJxlezJA86PMlonojMQdTMHeUIOqIedR8YWNC9rbn9nmVMR20sf
uALo8DyHtmstveCkphXVN+fM1h1fzy7u67BRYYFK+5p7YMFAPls/5hs4kudt8+Fu
QJb+MqRIF8A5j/YuIpCMXZjzXrKNuQ1TP+1z5sjM0Xe9z3aAlPRKoKFKGYxE4ylr
GC0s6Ng4wy7CNIRF4pXvDuRdJe7OclwZEabgLdH9/vh3PA6yJGn9UC0OF1xNLc5F
fGHZGevoli4DRv2gOpS0VHLIuFbsTIqPpDye35Nx/7eTvfcpmy8W0vmhOj/xXj+H
zS2WyjS9Wle/7jmHSiKek1t8zapdJotTJ/7TtgfEmOW1quZXnuxr2tSMc8ay8nby
+2LUpfcnTYT8Ao8poqQJ4ukQ41c4o3DVlh7R3zpfICw7zuIpwQWLm65AXDzmQA5J
Re1mdKDpPu/pAx/7ngpiWDlQZ/m2u+P4mUR0vOdvVKHS0x6LnPfF3tb3Ygs8sb/r
K++R9YP2l9dvpmL82nH0QMnHQ+/DAi+uaJJPEZNB1hxppVNI9qfP+UMl8zfCOQCI
LxikEFSqn4BIsDPUq0vXcpojbxKvDQOr9YOGidUm1ZysTvUuvtN5F4HQCtkIC15M
xncE5zy0ouXHxU0mXMEUuPgUy02YMxWquJexDOlId7R0WwzpKB9V2l5P873ljXmR
KMzIdhy98FuPicrbo7DBx72PeBkQvkvV8RQVbwJAt60jPxfRly9zKYKXsgkql7GP
th5Az7ZDq/MNJXeaps63x8To3k5TEJCVSQKifjm4QsmvM038VkPdL4MBm3HyVClT
LhyzAH80xSPjuGyKWIEedkdbtqpj8dcmzQGmphv29XluDQ4dM+aQdnYE5G/hinw1
27ohD52CrZkBbEUMnfTnxrRR+osEz5v669UTjBodEcBm3rNbg8vZ5v3npsnLNO5U
bc5qG4J+BNzDPZsuW0rYJOebWX4KQv4bbOcem3GU2pXYrcmEa/CMZ6wd/+GYsnI3
8qFh+Mvu2DzvVOMJ0BIF0aQXlhkhSvO/b1V5l05JBvCb4BBteyXnOnZhI5BrJTg2
z1VFa8UjkT6YJ31irHf2mNr3+7meQuocfRw4GsFor5p+IhB/karAYm1liJR7XHHg
11MHbpwGTJvfLaXM17hudmeNChyHfrs23M06HaaQhSokKfv1qqs8mBTRksL9qYf9
blnRQfiR7uYw5N4MdccdyPVsY1B0PJlXvzb1DsaYPB67TTFVSA0mhuoY/VkIopE8
nLjlmD0aMqfvlX6ooHniPlHXHX74DGb5wn1jnJnzOBGGA039j0CAIPuHONTqsApR
YXoclMxyRe85T7U1/DMpmU8hWeDW9eZWhQfQgV9IKIGDXNwA+MXi19vVkm/Mv63o
UDTWesCWSJVPAlTMEiYYuelwXzcfj2JDeOEipdnDuFJmLuX6xKtIwGecbn45ne2+
rlxcheMUzeC6I4FM/D6xktRHrrYRYtloQ600KqTGqNtyM8B6o18eSviF85QRE6Qb
GpzM2ooveGE4OSilxz3VsyZxmnHJt7W5I4wL/xUF2FVxNVfVePE7Bt307aW/bo+H
uMOvxkGU8NLYs66u4g3urAEGBWwZlf95n+WKOc9BttEMrlCcxAduh19Gqm7Avpeh
+LnepTTDLmrOMaOts3R3Pr2sVbZZo6PYEwnp9a4U+pmS1V3WQ3sgddg6xBW0ZjRp
l49LD9sfgBr9Ta3PuNTpVhrp0Da/6iHc+oeESKc1M6HiDjnSYHN+zn+bXGiLvdHy
S+SOHQceo+Bn+ZuMhomBxybjw/I/QMi4ws0AsKAPbZKlMqH6a/7Ax2HM7l5INCnG
Exw1/jHclfxDwJhIHoA5N3l8e5L/QB0ZIdobw3xTNvgV4aefg95u9jay9CiY20br
xB7AmMmFrx+2+vtLj2iXVMO+vW7yNzzcrHNt4FL8dnmX5/UlDDiqm7HWI8xul2q8
zUOy6SzpkDkFlgB1AwKodbBNZk/m4pzAGWRTGhNr/BUxscLloZtiTx0yYGaQT2/D
88ODwuTn615+TAQjbDP6jbNBGkd3i+gGYYqRC7GSJwDaKQSrUPvUPZk47emMvtxY
+vd64wL2VG4GmTaIBCgTgqVKp9duNLyKjm4zg2xY04ds50IQQrq+DgSOg8nJ1ji0
WpbQKzTZysP/HlG5YlQAnKICYC8f3Kia1Nip3fyj5UMOUgJk1R6iZFH5Zdd+Soaz
noryH0htAl00OXQ7RNHfyBJ5+7NYZ/8kkRlc+YNRkyrRcgPSeExqlQ5XlXGqOplf
LgMj8oMDVxp/arGN9m/h3Q0/egGNG+jiNqrUtmupVJHEBudp0mD5zpYtwCNVGKZE
gcMCzuQBdnnLOI3CpF0mHohPkW56/8Mk9e0dpLQwIMttSd4wrKe9VdQxiLjG+out
K4u39/yjMmERCfN8TSPkMmCHuppJJ/4Zge9Nd7ujXEYHt44BXkpMt6wXwM/WeYZ+
1i7+6tc+L15DcvsI9VhMtI2c0jBYlhxW8iVzbF8Gd/g1LO1uN4TKkT8koSj/SL+q
5cbGknW+8+bhQhYU1Pm0gfi0j3R8lIxuFQDe0720Q/cnwBmpLxvqZzT7PEhfUMHW
0Q8pFGU1xlwdF4SYjQPJlYfYR42IL0W18dGzPMJv4P//d+oMwlgTCWmE/OMXbi7R
nUnu4X13t3N4WDblexv7lsZLBuem2U4ZRGhDhZNmlcOWd622dg6TO+kbFkpSYW38
5lgXwx0A4Hxsn02Xy8FOQb44b8CkETx9GtbkQzVQdsICO3bCeKhrcev9yKTHE6/U
WvWxSG05G5etDO/C2HdIPSyGetevzMukltGgzCdFf95uu6HkTPYNTVGD1PIg4A+O
H9haTaS832IUyQbgTVCeeP+qnI37GqaVpkW99T0pV/7i8VSiWY6D2Iq8f5issFYU
70e7vv38P690f3BfPHQdfxDiVscRycNTVepRARnLhtZnClscH3gN1+axrH/o1F5W
kpLkhWFZMZNm5Y94gyR3r0fymlX2RTBRt4MVGuf99zdJcHJMGmXShNOXUDNmsnnY
xINT/PKwl3gxVALgrmjdAHuwSKzbD3ZXAKob/68fhFSWPDwc9khlFsc0AzCLE1Xg
B7JAl2QK0CjMOsn9276yzSfmZzrXP857oihY0cwxNjsQmMbVtwWYYtewuxHIAuRX
BpSWsS7yOZbwMnRpUWhtcV//TwYsQ3d1LDuegvmLXo/6xZ8NZT6ckgjiwEbsMfuh
29JAejCrLy+DMXvWJYVj7sfjWKRp/bPY5vKGNFVhPR9Ix81YzR6g2+Wrky1jzO6o
PzFaNjeJppaI/vEZMUaHUA34zEDg39KVyACbbOMK+PB1SWZgKeTXjXLhxHxIv2IF
sayC7tvZbloWdSwwEjOqEBTzoTZGI3Z1m7UqRohZA00pys/HRRMtXfA3FEkjBdQT
sFxX+WvxuvgIexqLqnlqZmwXfvwtH4oEjJIJ3ZOstypqyvJ6hLq7dsOnJUJorAdj
qUeDYaYg2TptRyytRtoiCB71EArcJHG/0zGWmuHBYufO255NWlNs1PuXTIAgsqKM
kUNsFDOfKvNz72Z0lu5qG5wnQYj6dRjWaJvXk5XH8DHZHQh8RXf3J4qszsFbr+lu
Jfx+4/l5tTs7Hcsl8SCn9oxAXlltvxIGLeVlWwEb5iyTeQYe8Ys4GgQjGqX/Ld9b
m4eTmEqHRA/ikKY6uvcxdSI6JF44wPsLXsPnjHUTpad8/fE4A87DKfxvg3g+oTnq
nOg9KeAQ6CLK3Jh+5f9TX3u5+DtJasXjpZmjMXi5cUZ7tb9V7NCh6uVZzX/ihklI
1T/m6AEToPmU62r7pbgkJ6NDYgYFssSWZIRAL3my/eVTNUz+O6+1S7BhJQrLe1wP
af0F8jnm8NeshstsxVyxyqSVpB7mz20k8JBdagCxhyyZ1GmRTyjc0kILhDgYozDR
+pixGI+FWN5zHZNmexhtgO+dlXEJbqW5vawexp/BjzBKRo6951BAFl36aXELa0Q9
nq2xHHSBEXzu7f1wCY6WTjEsC7c2+6aeqex07+dCcwlc0dAoBKb1num0y6ffvoGV
h5McjhczD2gANCUXwtb1Y8KXBvy50tEA118HZcIArizaJ/YJuuD8GawOC7AaMWW1
l/Vhb5DPKBceifNegjiogwj2+/Lbqxo1veiKOY3Co7Gag+r8ljIcCPIc8k+UfEpU
qkkr00FdToT3h09rcwwpMh/6WLteCm3gWLzDoSw4yrMPWSzz2BBKzMI2t0vnw7b3
rHTnTIH7W3apw9orn8nPzxc4SpK0XgQuOd3V3hZma0MVKFZOJ+Ii4kXFOubYTvYH
TouakIySMf/k87q5zCGUKOVjxJciBwPJqAwvgKCgahCvjbOVFDvn3ul7QqVA7eTt
GK96OXk+hHfGiR3GqROxtbZqPla0vuLx78QNMoCKZbiiUn0J9nsW9qcAugOZvY8o
335s/GEPlm1tYmFzR73g5VmZOR8cqyN2iVsSVJbqNLVkR6YC913RYBaGNbIkwosM
0zRtm8WNHVytywNFrskPy0X1GSUEKO0IFTGwSOOuFWHKq18WJ6hDjhu4Q0ZLN4B1
csjuAFZLApxHpF0nxzp5L7s7F0BPDMQ2XwhyaEcwfOdhJSqs8C1p9GBQ+MFzuyMD
8tu+Xf6KQHPVpEoyjx2FF4ZzY9gDjwj8bX6x9/tgy6h2X+Fd8GCMn4T9bxrJ+GFC
sW1l/WkD8afJpK6iwDaHBYbNYhiXGieHjXrxN1wXxvQ92XjMzmfL5PKI8Db7IjDX
rrer+lHHVcp2uYli/Qu6ZwTsV0GfHDTVcSwk73pwSU0ap4FVY2QqOmgn74Kvox4+
8/UPSkmBYGd1EoYrC20obyzZV+zddqDb81bZGkPDHQeYeA9pnd3anVVwYp/HRgrO
3gsbD4y3sp2pxaVlfnIkC46Ne7XW3He64b0p+uqIoaE30jSQKNawMMNxRXNCjBTY
N1wyhuSqmMfI2nIPKvVCoC0k8tq5czHJVW3m+uKMwPkhxtTU5D3LNmqC8JoVcaQk
5ROEuhqwvsd+rXfEE0DFN8auwY9H4r/kbrBXwylFUmw13gWNBATjCXgB6q1hxpbM
wTOBjiVAuyp0c4IReCaxMNxZq0jVXhtqfJ/tlFIrz1N6xt2M0nMc5gGTKgaTTZmk
OQ2gu5qulaaVaOWboGAiCl+t5r671WYz3ZkX8ddpyeW2XdwBTb38HxKctMBVEDf7
zHg2u8DRJiSJUmY3OJcer+EOoFWoRC6u5MiFr1fqaBu0OtdJBHYoAUbunBif/Re/
7ynDzVUnjxc7eh+Yc++obk1O0aZuh6K4SD4WQBASvG5Cn+a0OM8C2kZY0xnbdO3H
SWLDQSHqfoLFBuUhbc/VeCyILXr/zjhnmFWZsgb/4mxQcO0Zh+aHJuL8JyU9Hgvo
Nv4NRyOslK1JiUe43A6WbOUr1rHwS5OCRQHRaUy31x1EVur5OdNgWSwR4eY/kTq6
KOLTBGALHDBLk92+b2P3iJdZqnBc7x+bcOuAHWUSfjFS94ODDBpadP7zr/6arrV0
CBf0VtK6LlEyHzfbBKhuWVv96Jb54ZS8dR6Wlg6otI9LtzbFhM/TngOxS/i4J7Eg
Q9iTrZ25OlT+3TSpKkBlxOVUNuac6SgqpyNHLZQh+PLy/kC0PUYUWZG7qllRTO4u
o5ZkJ0amArl9c0IgVcReLGJFaH9q8kBVlOYSMrMtdM3ak1yuCUhn5MtEKPfwYpr9
xnKQ3OUwBnw/mRJSpBPzzhOwb4Rrj58Gg8GRCqK4DUsU7d+oRCqS2ZFrFMsXlwgp
zZ3v7jETe1xES+GR4D4OMokRwrS7PC1oAJKHq8+uH265/jnultkISyCOU7nwpBFb
KtZr6gA4J/gAQt68FoJLmT00+Ikom0iwvzOGsLvIcdDswBesXiWAEUGIAfJpCL7T
SUfbgIBBoIBEdLP1kvd/RWK9Z8eSJvRNUn5A0ZueiKJeNyD6FQTTkXhmlsLo3d5H
uXiMaH5OVZOidY4AWy86k6S/Ruku0gGkKzqL2XvqwF2BIktRohX81mp7p9HRLClU
QIWdhgPJhs5w2DJduRfYXYl/m5JFhjcwyvgm+0FAH0Fsb6P+vzacfGMNwbUondCv
9g5tFCO7GZr2XO0tZqXrOLJH4F60DEIiNxwua5MAXEKPOCY1rRDnxUp8peRy4T3O
P41KMCVx+Za0Yla0jSnWUql5jBypIYNJY6LY1v9spmV3wQhxkMw7fTeIAyEblGgg
7R9pvrer/iOBkoBDZ4H0IbRsjEKJJC68tL9RI4fIEawp1gTfHguyr9/nEvgoPT4W
pwk4St2BghcZg3/tMTKFPTUZDyGYkt0auJN80xE/SfervOp+qPVLXW9mfqiZIULy
HufowWbHezXVOlaoAj3A9Ug+65uuB1o0G8Kr+pVpbf0jEwC+XN2z0/gmsmy+Wxhs
PtRHnVYhPbJDUwH2Ks6R4FxYf5Y/lNoEZBlCssGuAqw73B0/mDyuzimznx3P0ajo
nDu3DuDJtOYm/Z5dSNGDJNehY1wSfhzZoY4bHMMi4NYefTrvsx3e1Sk1NgqsThRt
9fHFjzKLflZ6strp10jPL2lQmBDnry9vP8aUyIx6zU8McWQRH8Usqr3ePWi2ns8J
2rY9KJu7u/nCv0LCF9r/EGQ0ItTHErUivcMfGmoLC6eg5FjptL0UsdPrZYwpnVxF
nCahPiYaX1cLRdL3ir32ikY2DUj0clxYACcx0729raC1zyL+b6GVPFo6pohZ2Ljx
iZBtCon3oLRxPH5uKKiGVvFGfz/iL7pC0WurjTl/vIiRKJXWms4N/Wnyul/FjSjC
ezciiCvhBctRvlintCVD3ErU04Fsr9nt18AiV8535L5kt2T2xMIsTcb1xfwxAd3a
ZDlA7gTFsQ5d9atXzCwab/R7T7WS7FPu55m8bj2Xr5MgrEoOXGwreEDkWFSJ9726
EEMlsFxdm+cLEId38X38sZmxADdH5ApwQEi6EcCEX/tOhxyf7xjvZvl30nEMJdjJ
RdWcKakKjBy1avjGvEem8UD3JaTlMDG0k23QXb/H+r96zbIZwXLkbJ8+lTP4KENd
6YLUOmX1VBxBzSV9BbLBnQlh/5oZ+/rBIGWMBp3oTQ1FnWUDZwj2hzE/Je+HxvbB
SVkE4G/O0ywJkqOKqJXsOhiqo9rW68Dhwb3hjDYa//gqvPKEJQsdoxNQz/dmNEor
8D2voFVS8Ta9oRC0Ot0DTB0jCXaLDeVIuw3hvpK5pOKGjccKpsi4oFeWmTKazLPw
S243ol5+UcAvsrQvBC1ePCfyWT3zOWZN5H3/XFrufrgMsqR8NOhaKt4M/VGFU0IF
TnI+6XE+peXVPd8MoYCRxQGb8xpVYXM2+WJLZN8BBzaK1+WuiuKuKofPeN5iG0V0
Ix3TrRB6sBSkqYiQ/3WZ8X7jasZ9J520q/r+q5/EqOMUGrrTkhk/8QeA7nq9DU5R
FS/I08ln/1ZF4WgmJitRceda9HilqMzF4XJTl5Jqi5YH1k5n9EwxyhtP+9L4B0m8
WxKPDX+syNOI6btkH2KrOF0YT3A8aDi/SQVHxnqAJFPH1TOdpeqZT+Pzx4djt1ew
fdJY1IScJJl1rUWGzWNxa4yUvcOEinwCUbAfFfh7sP2OVrD567XNeHgTGFd+a0NW
cF7AaKxXKGtVqck8Gmerms8Hbpjx+tu3s2qgTzX3ivAffEsrJRNHRabQ1Yhk4vLv
917jSxN5KzDKywGukX3TP2pMecyqda8dgGyzv5QPsCupzs3X2FwAngPvgnP6aoM5
Yl/Y9FaocIDelY+asS87e7s4CzVEc5SnNJZs7pdTuApzVhS5aP3pHbQ6gKWid/9a
nKsumd9hg8sqRVjX2EsRVgXv0scC0axxNSQDXolrxwjN8ny2d9nmEOd3TDl9EuFk
OqJitQoO/7EbuL8R4ewpEOEnSzcwzTX20AmobqftONgUetZMJkZbTJYTZH+gnPX1
f2dODHtfwXeS81t3Kau7gvilsmPU2wgkX24yR7tpvCGNBlFQT3yv8C2oAWjpw7Hc
iUKb8B+m/x0tQ4B4wgxJb9wTF0iRST5QOyiz/Ag2a0lEfrfEd3YbbH14TtstH8AG
kje1jsLvvZ0/6QePhpfW9dKh9rJHLBGjND8Hgievf6RmaF6Elu6+t1evbHnaEw3s
SG+WQCMnd2K+lJj7R7uomlEuyvSdMt/e208E0q8l3iF3mE58liy5hYDNnDprPcCw
XEdZ3T2J495mQB0BO0JFCW8fC/c6KJ6xztGWvSshwHeW+Vak5TZNVqwjGZWLwymv
cmgtBhQonkoQSchBkGCd83Fte/mduC+YHo6uwiXjLGUGz7+f9FgVP1c5Drs8Xk7r
LS1ZnLJQN1iYIMTTC7ryfWVEnmyjle7pJecbgjP/RZMwnxyjIv9DP1S/9M/MOSZD
n+XnJDOUz6p53XhPK15qVYTmsSqvIxBM/Eu2xrknCo+BgGA590kcouTMW+qe1hXq
oa4EeqE7HLc5tC2jhVTMzVZSwMaI3gvrLq2NEhkTIxk6aMtT9nqQ/S2TJ4Kg2bOw
OxG5h8WLNfUf3CtfK3xJBHH+rZV2vVPqXVxHaHXz8kG2r1MQRJj3g0V87O2thC/Z
SRb//OzCEjWs2AYbtEbp0ABUHp+gFJSPWRWmSz0nzM3uMZ09ZP715t4SEuFn+naK
8W8sDIiIuW0vqn3LN5EdE1s77I5ExiBQleDcurPLpgfb2I793U4DDOkE4kZWs6jq
kZL4FL8SMuF7r3XtEnTdYo1g1hCWxSuxJlagygDJQJSg4pvp2ZmTHGKJCkYoO9PF
2gxhbQRnGSZxaRgRADV2J5AdFP3lRom59eD5zAN9A2CqDHr0ay8212aCrg/r11xV
qh3dBuZM33F4hadhMv8OG/qJhgkf33WDbv47y6fPfyQXx6lDv4bnehf05UE6LqSm
QfYTRK92sZAnpTrQGilrOWTLW3Mi2EmmO/e573b2ObG8foKU3M/+N1kBcyBr/Xg6
MMAtQAGIoDGmC/E0LHNwdXlfZBEPE6MuriycyjLyYgr7ywboXoUJb1bCVv9vOKaL
/QpX2R/P52hXiGLjevzbFh/l5AzUDx0Q3hydYdzi+PtieG5QXxPzjUczZMken3xz
zloEd7r3DMuMA4IzN8dmFUUqLJOlBeCjI/m1HwewvpdWzwwc2KEPHQR5ChDSzug5
oY+eOZovidy4LLYOmLjxtZ2C3kq10z6ReR04UBVPQbGpulXYG/Ao5LrXIuTSBluB
+pUOnEFe5Cvj3qWa5zsYembcTzNHa9Vq1+GkqgSrAo5tgbm5Kn5bs7DLxjX0m/3R
qZS9pfkIWibG1gEj+neRuJGiisFwrPV708xjo4TlPFt/Ptk/+Fo63Uq32J1kBYP5
WzAGFuSPxykd3AamDbJo4NE41k0HZ13Gx3BmtuXALxpEO+93RJy09h7S3i26I/r6
pxYVQ0Ryt1ul5qHyskwDpXeYqF1AcakvPlG4jAPoya8Nea64GvpqeSA4OnSpcwCN
Zozi5rmeCF3AHny/TCiP6dpn1/Pc5gQ8P/DO7idoSlapyVvrgDg0/hXM+njGanPy
j+rPPqz08A+P/zs3+D73TLxkl8tPho/STeHLNtNsMhZfgV40fDQgpTrrRwlhCUTy
u1YbG+1oyjWsypeiM+3iCoODADggNrNtz8qhYiyzQ27WUjxx8rplPILBAouGxWBS
3vDvf2vJDub0UhCaZBh0rbvV1BBUJ6KbmdAZIQrrL4oN32NAcCKEMBM+O6qAdDG8
5CdkW3Appgl0c/ADZSpyFcCmzO+P44DlJC+eK52Jx+XR3hmR6UE/I3UZpHbKgCyL
5MxR7NydcMnbTd6wgOiixYabNQLANgcBvqGSBHUmY0EB4QTZfxorjiemU3vfZ6Nm
av8GoRH2Sq/YtSro1Ql4Zg7XPBK5aMZV7HeiEdTB/KX5RNXJCr37I9SeONWMxjHn
D3TPyuaF7OT2zeRMU+nZ/wa+AsLV+W9XvIMdASe/KRI9yTpsGWnSroQcQZOy4MQQ
+NTO7BHeQbN027lIoUc3Ap/FPdYQPmEFfXHRpfq9dBReu1q2By7eJxXEu/VPB7A0
7Jwi9T5g93o3/U/hndWGqru+uZsNhH+cvXwCVdSJYG8VvqmhLi02xNnVOrBlNQKF
QhL9wboTXMhnZagZi4s6FXgCSRwxIxxQifIqRpn1pzx0F/ecH9XeaUnU22BR1JkA
MnbP1eQvSkGGIoWD+od9NG2zbyYmjoJmg0uCg6LkLJCO2Do5Hq/oblAGX2Csy8il
F+Pad5wDcp5IMkXWDhphqgYw2zRU1JWds3xGjEI2fXO0MrjVaCxIRPq//X1i51kH
MAhJH7j4SDtBZgK3mwasreJJy4NKHwYbaw9PEQkUQQFRghglUCIDnhogrXvWYHLC
0N/+rxpPiJmTUyumYa5VUpyA5oQZHqovjXYA8bBPitnMeZgSCR9Fo1hhG1p8mnrJ
I3rj9TFAZs6QNHzTI1WcWYkLuohcYUmpRLz3wdoBXWEwxguUGLqOpmMVybQi+71C
bf3gl2E2G5CdWoW+bHVmRBBM2z1ZQLLppLSd1jYQIE6nhi7HtZOptG90TMFtypiA
c3rP/h3nBknUVuknrhUhBSHREmQ/ayb+VO9pxyqRSHHmOJBpH4EgxpwSdXnkDoGa
bEEXFjt7xtKXgHZ5JSPQhr5Riv1Q+U2/BwjHmWYPtsVGIFQTtBdsCrXxU65No7/R
IReALonmaii1JXZlXY4EbO6re3D4f0axmJtmM8HeCqQka/5VcHgQigGnLDB+G/Xv
Sw3taWOmeuX9EMGuUVHQ1n9BN2YAgYt0HD7w0GQ75J/mrJ1u8JBfix/NoGEbL3Yv
HLnRyV7j8eNrTKxRrwOo0BO0wxBjsuKN42kMG6YZx4m3+Cdw0RbQn03sAKT/EJTs
PerkaOD/l6BuAFPSb9oLxBEBt7oAYE8jZ2MsNks05TiUj0QDi0DhSxdd/LjqYWi9
MoazbeA22T6wCeCrh6zsFDp07F3S/rg+0FhySWN9/l7Ep/hgEVQH0hv0JGC+2Sva
UZzcmpqZXul1fs0qNhNolV0HzVsnsdtSebjSx1WXQaRrUxjYOnbkuzK9oCgrgiut
X+ezpgCeCIDbkUZmHlQDItnBHbzDGDZ0TFO2ap8i1vzr0qoD1Kf7CnSw9cJt616Y
orMtax8VK2IKlTMmZmyy1Kg7hyyhnzj+v3vVgKxiVbCp/IOcEE4m7ehK1rat7jAW
BpoFrXfOeQTIbVDDMMxSOiW4qN9nzuhhtWwYFx3sSA+4YfUuzWA+tW9Bs9HbAlh1
50JhSSsKhn6UePKlcI2o0PAdo1R2+uJyKe6J6I6y/9oH2G/y/0+X238ehg/kWgAc
GJ/3imQLm4licx1I3cW5K4WS+vOk/bXKLJouJimrtwlmO/XHyzDzg7gDDPPFZRq0
smXNaTi4OxgWopRL1KvUifd2DW2D4vNZtG83TOnKPUvjXAhpSvDHCnO7bLJMKjs6
sOCXQo1Lihw1yHklT/dIAVsf4x/0LWn8GM6bQDI+ATvrqPv3a1dTlDGTDGGMxnSb
OqKBaink4/OJGt4WtzgJQLIOy5fowXLp3rHFOeQeyQwHTOi/krQHXn23nSIIV6MD
wTi+hw0tCpYkGRTkYGbtmy9nYx5T7PEFiw5sp5fUXPo8z/UjvNlzqoicNc7LTeXK
PWTcr3BygzJcHG3xWm7fe3gwe5/ZryDYjCrTx592tSpUGyX3JcUSrYcxvngwyKdy
lElWHQZ4muES7dUth1PUFZSivJogG4WQfSy5hW3VTFEaIo/k9iy5JPhvmTjcA1ze
BXZ8UpxU1RrJ0m++vfhT2bBEVCRf196/KFsnro33y8le2flK/q9E5QkZGWpTPGes
SUq2oyvsYuw0HLl+ac6ZiGMQeEUY9yOiKILvPaXDGkFYi3tqe20qPB5NV2Kk5s6B
8ETwnJ8p0SpFRAhcu1125zOxgKCcqLOaRWHzHpNW7QiMXJEpXmpF4b422MUp59lp
WgOMSPiOZoEvHaAQFfeYnRixrd7TzxSGZRES7H+lEXb64WadCOagn4LrjmNxugwP
699qQyBFYFQ8XV1Tk/GSZgIQ1SlWLl5eccZ4zX5ShuCptr7MOceN7zKmhsENEyPE
KV4JPsi0sJ8Q9pFDRR2ZyMvrEeoWzE8s32mrZphaMRceJ1E9qQbqPUF8rrlV0Nbm
yFndVmQ675gGK6bImfgIzAv+oTtI2FJv9nA1d9yK/eRkgo34T/aKnGZZ37GfbPnR
xVjs9oGc8xQaky8BNub4rQYiiLNq000ks/lJ5SdD/oGDL6PlU+lXGku/5w5MoVuN
qgaZniDSmbT5KAqix/bc2YVGkI2IL3C+vKCx+Wmcpto5cyYgVm+SpijhbhwUeZfa
+pyMNGiH/NUPpYS8QJzrKFMeU+y5BhjIltH+vjIYDipA95RILoIkcPnR+E5InqpB
H2CDeHnVtrqskygeKDRaIL2YIEAOoW185+xTLbn8HcCWC096n6t4kad8No/hfvm8
aui1OukTiYtGdheQddq8jHaFYAyTXDwVFVFUdENRyuXzx0HKYGXAt2rw3uedzPan
1gltJfbHUHs07hzxNjV0QIYDJjAFfmlPDyR+/wQBidQBqy0oxlqLVM/k7OyyLLdY
NIm6++sv0BNSn4mtSDsVakVQKvcw3QheZ15obLJ4LSjGbLJ3KJYLG52f8czRn8Ck
2MOZYIegGKkRPOcsjdw9PgHMbiAtD9fKglrxfUlZuTXt0S25D0rOEoNJV6jmk9CY
/Ujt02o+xsuUhsAF4SVMXZajUNL7rAwXh71t9YhWaupP/cG33qnjyicy8iexGw8B
Pgc+/Da8QRDLpFjxdq3ruxl6+4H2b23ONhKU835O4Enb1M6FLPKWyOtyIkfxRyok
HkBD3b8CQU1kdNOoNhr+6deN/DjNBbvx7u78NapGSe0vqg4i7aSAaC3Qspl0I+I8
cYSNubKCiTwHtV8kbybv04qhiF+1LPBtC+3eCYFz41UToL7T2BVtBA2GJrw5rc+M
dKS4+uqviqLETCpTV/SekkMYx6k9LqmXUubrgp6VHuoFJEcueAv1X/89yHjncK7H
tz00mG+OkGgRzBCPzQtnsrQAJHEv5wipSpCTOL/M8Xi/hxL3WRC+qK8k6OZzcaTl
NDd26cNnKCj/TTP+ba0IDeuu8081IcvdqtJ8cj3OAdpmGbG3h7UGlUArp+DaWll6
FiU6PU0ZOtjfxnM85ID/V46ymtYleTaANl+6yYvf6Kbo1KwERuc0uzz4GSxLckU8
J/wU2uv4SiOZ2eOFXDQIEFEa1GCCkM35v2BLu5W7aMF7WPdGi0Agv9t7pJ2ixFf/
rFH0M2R4nUUx+ACgGVw/zPd/iA7FwwH6GBWtBxOZEzlULtcI9kRaJi0iCfTzVEGY
I0sDckjrvv8AaDWUTnQQrA2Y2CaiGlRD2bacOywOgs3El+ZM/xFaehR8WVsdnPCg
ghgXCMzYP+xB/1jJTIytJhijXCH5xFU8hWrr7HfqWRgaSzRZQkWtoc8zsqAFgGQz
Y9r4Y7HGySd4WLmGn79nCrc7UQW5Ieq8CG5oOUWluCVCj6AEgPB0yU4NHHEaEyuq
Q2dxhz5qeTBngxANlFjSGn3B31mb8EElUaqkW2ozOdE2aAlkxOvfx7nj6AEI4eCC
+zq+mGDsMiBxWucmpyB7pcZBGa/b0GR8tH5bNj3Uo3j6ZlSnIEr6A03ynRvcBbF4
o6mHvzK1I+n2t2l7n3mxdAWCFEj9qLcZm89Gj9hwYAa/JAieJdIEoDqHfJL2DNUG
4pqsAPi84arqqmVHYnCj2QewUOZCECzOcaojpSl7fqE1yq1v1Gb5GrliLrCfQoVu
cqjxvp5TZiKbd9tAckgNZeNIK5mMmCRopxyyx4iKkve1db8ECrbSk+CbpeuDQ1jv
0ReyLW+ZPi4einXJl1xPVI/KjSorNOdtQLQgfZpJFEke1zlpeQdhJeGITFqMixal
dqIDCkFgEAxzhWidiDqFVWaLNPXvedJozCT6/RFWjQI56mr6lXbw9p5bX4RQXn+h
98RFolLHg83+Y2b/cyyDMgl2vJOlZZl796Ue9aE59FeN1pRQzZKjx2dP2+b7Y0i2
9ywdoYS1doGQIXRJODSsQt5kKin5X0qPu+40KaDQP2VU2OmyVWfuVI2MbzTwHEtR
h/Ujs2YzFY5msVT+xnneRil7SxrkixDUo0cdoo3SX7SAkrRPXCxBSSO5Es9wkpFQ
9wNg3nfzrBodupaIWUjzNTKAp9lGskjZCKiL2B41dI6eKVEXpZMWEpDDfHU7rPNQ
4/bSqsiiTRVeoY662A/ly/XD/NFvmwvg/yMyBsLcbJBPASgpCZxYYKdBD1o4HsZA
AhnBhrPzmPunf+PsWVuRa/EBXfVRX7ddsVFjPcpIMPfHUaQ6ubKIlI74okNdwJ7K
2nAsT+O/5yi+1SZ5hhcGL2LYd1SlmuEaWrOaSUIc6jtB58WSEg6ZhDkBOpR50bNN
4EaTJqUhuJ4vmuJOOPMkg9qhdFFLSdpjs0n7YbciZgQNZGwV7NRgVc7NeuGai/Uf
oQpo38pwZiD1WWC1NoW1zMu1ETaiNtUSJx0xEX8WVMALlWOOm5lONSDc0AdyJWtP
DxtJS30IZjK9GLk9s4uq+aOFvdUnL7I9Xk8uAae4ygFrtFYgmhmt+jiIfQPClVMR
UFO6kG1VG6a69OX4Sn8Y/GmunFR7glP+IBoiqCPIlVzmbrjwXc4JPc3W2JUPgCoW
shQ+0w8Ixl/Z8kuxwNJ8DohGJQqyScTrnWym66reYo4hjhHhzJdfUR8Y2Firr7TL
kFejxSZR9MQxl4Vfp8UTyYpSAKIqmlTANXt+ZiswsgfpQOrIv+8NwNT5xLWkgs2g
ObMbuA2pfNbpcnsCLgsh810UwCV8xBBpXxZSGxK8AGBy4LeZ2kW/Chb9OLiDHvHR
0PDP5drimDDvNJutpZtZtd6rkP/9dY0NpfKIJl4lrxGATorJSTEzCGshKC1/zvJ0
ysF2LmJbieMzgPPzOTDriGcS7uFDpTqTsN+TvWubDFTdVWbulqRGOx+NOvmvKmDj
94UkKesgnFKN0IAMmT6Q5hbpB1t6r2IkY9PYkddaZqvAfF2S9h06vTIXWrAWOB1/
P2DAPv4k76XrXui7AWRe25bxhiIzBODQUiCsLd9JqLdQtehebo/4Rsbg2OF3I67j
K+DOXsRHICr01v0gojFnlw/5vilcL10ozjbMi3QNRrubtW9cgN+/avC/JZLzg/wW
DrJ131m+uSQC+JSC6NtavK+eJ6peu6rd18zjtTNH1js+Z4u9Joa7FVlJSl0RVKNI
h+hauplDstGYPhD9i/fUM+8y4la0K3mhdQ566yTcgjnC2P+oyn111Jz8R+JnIlIH
xdFBTjwkY+SEioA6cZxBsZoRu75YBgNCAUuF6SsIGlMMnMRBsygr5LA3FHNPk+1f
UPYQ0YQSgBx7onblW+ac6MgOFWfA4SprwZsdmPrD8EwWOkoWsAGbjeWDzPuGTdfO
XMLtQpFJjQ6AQdyAgerSyAoULz2LtgL3WSLcXVt+n+RqKTUoEiYghJF20EYC5aQJ
iKV8Awuz7ELGEwQnBFo+fSihXMHOHkuKpWDntr3jZ6N/07WGhZacG4cy1sKh9CIo
YF5c7klHQg4wJgkS/h02e1etSRcuJCq0i5LcqM8DNG42p/AU/34asBQiDV1q3nea
+w6rLK/gjxUOSDMqUsVRC1vlXooV4DzjwGaeN6mylMUngLrBTMr9m5F/uZUUhWeL
geqZwQhcQMz7b28/r6tV2eMU5nAX/atH5EQ7TvYo2oOARn/V8nH4u5RRQhozirnR
ksqoCIR4jnx6Pqykfz7e9JMF/SPCAsecLjjv6rvB5m/+41hfrOZ4dlHDmnl0psdD
bGsiCyJS2DxxfxAEokw2M56yupyrQEKeiF+yKWcLThsOkj1gWXwSPts+8o6TM2oC
SOz9Yw8QYDJb9Kw4OtLsxWzat1aburkjpbkse4nna4FmX3sZot7B6GOjd9K91Sbk
h7Y2vBNOdxJSGz+nTZyyCjNzMXaYvq2SNGt1cRnm6ZCbKtYRFHh/1VZQugvbJ0ZJ
MVQrHvAdIPhuJVerlTvSZzVytJ0zqG6Nd7JInLptHCUUBIOMdKz3AB5HxNj3zC+2
j3299X7MI1ZysDeFsgMcyll3eqaC0povQ628oiDxpsPNoIKHl5VQznI7bUsUyenq
BucHyT21aWVZyBWREyq956s83o7MzNzwhlfPPhgxOeN8GpgMFPKIIpquQCwpX5P0
xL8kR2DtXs4JcqB4V0MH1n5X3gnTI/GupeFD0xeM2Di8o14wEb6YmL2VrrpSwIGy
FlSLwnf56ghjvhBEFk0wdQgJx9Pc/PlDgNrvuMZ5KtUJs8xQCQl3HXt1Eyqi6H1i
2snXPoskEO/Ns0UhIAJnsVS5Q41WcZpPshu77e/ZxzAxui5cQFH9NVbALZCtalww
Vpy3qv6DC05nvWceyUCBpsS75c2JftnwCrSVch8r2Tj1WzlX4vWhPcgUpuJY7+7m
2k+LFXB9BrD8I5YAPoZQnu81/+9YeAgtr/Qk3BsLWOnvdBqrcZ0iIFvmxS4RkC5O
U1ODPG09rx+WIERn40KQincM48zCPJ1Ss2sdjxHqlYCsFtzpnLZq04MUeSry/fWF
ps6ctQ4rBtfu3NqrcpqGztuP9wsGlYfrnPJ4Xc/wAPp2jRwADS95xZ+eLN4e7vuG
BIWDq+efV2LOSxxZrzVmw+GZ0iBuSjIunEA5EUslRcRIOxyOI/eALjZzooflsVE6
8VdLMzPb3FHg7kpJKDtFCzyarvcHViB5iXDEN3DfLqo6NarsVzupAEbZGWPTxFTB
ZC2GHsgVe1i/NQpseFhzcXiy1foe3olAF7TgSfUTsuH1DOwFmL/gt82BnbkPtAyv
TXo9tpc5jmwHO83h8pagFvP05lEZ5498tMWHSXkg5cW9/Zv+PdSHfqlpxDEUNfhO
YdcPtRHSq7aphpLDO827X7ndR198XQ8+nbf0V5UpO08fSaU08rVUwUiuertDEeqK
2QikcFY/dRG+6QdwNxSaPUFCFH6AO0bkeGBK2ij59eZ9p2VSsGELn3xdz5gdxT1q
9vBMnx/qxl/n68VJdbVqGBrG/IX0T5A1J5TACettjCWVfDEQWxbYUn142tyvf4HS
wc/h3R4EpBcEZeXxu5eWmMyy4SstztywLMmfykC/eT6PyDCSS1jBvuNvwRLmfV2E
JcBmbd1OVfTbHpccMYtIqb70fevgmDD0L5dQmyZqCIj4INBBMf4tOGBJL/tODDsE
DwZoc7Fg2BvL1vFbSLjgcpBJvbI5DsmOyRqPA6m3xQ5ATVygE3TV225UMdOKwy+l
rUZwMvPZTKcsP6spZjTP6vUfunnPqwXAVHnxI2PHvbzZYv2u5aRSHJXhN2nh03Kn
3TsrQEGf+teIZTPgEwpSlPV1GIqwHBw9BwxEV4rMPx93ExcxoC0ckcsTfrNE/+fE
Cqj8tHHL3eTg4VrNjPe0il5aUrRC+03lkvfpuof/KTmXvaTMOcSYYBMznabzlktS
Rr49/4w7wx8lB6VDbX1hpQtAFNOjvoxjdtPzATvn4Bx2NECIOMofol6ma8Hu65/n
kvhQhCM2s4OlXyIVq2eXNAspObihCAFhii38IeK40qyNjsFx/dZCaZ3YS3qOtQvj
BhrA9HiE8SzpRLz927N7XDxx+Q5K5I5+5JfaezND7VEmqXrtYCXG2WHRqU5YSvT0
bt7spvS3ZpfBAXFQfxbpFVATWx1ht9RPsRM508qrIWNXpEmc3J6gd8RA9d5IAkvM
WbgOnztaR9JBBJ/K4U+1FDWYcsOr6QtOrriGQY85veIkZWgWQZhsLDJFnKkn6TSV
0UHAA8Tj/yQdTB6UrlFu7phvVE+I+a+Sjk8qyIRDiyhli8mF0gNNu+JeQ8mq8Q8w
w5+z2PUHeH/NrL8xIw3MRcjcJPO/b7Pt+VcBWdm+gvMSu8GexHB7p6VjTY8616E8
oCVOTR2ilQ4298/YjsMmUC3xt9PMWO80kiXBLsqg1skY/XBbXLgLHuEMiB54DIli
XUohZhLskA690m6VGKY3O2HYgUTk9dNPY9phT6WA3rebrzNQZAo0LBl223HxzpZn
V7HSva//5OtN9leVZvMx8q6Xp9nXUpkIsCFiS82i01HWweFqduC1mBhcJzImm0AU
XW323D+sGP13tZboJ1C66a2cyMY3gh0ikNyips3OX/DNR+VN1GDCbYKO9qRTXRQo
1Ld00VMSesew9FKnjMCCF6gvOhSWCrD4orFsxQuXLFunqwc6O1wEijQpQa/6tp0b
FGAMCFJBVSZ+frldLaULnWxbgXpJ8MiIEmdDwz93m+WsgjlD13oekRX9/5yQK6t1
w4krzCLPrJRBUXGvnnLUGQBuDzSUep25jJgDQJchNool8YbYI6BweSpw66bc3wfA
s3KvJKTi9JArm1z11buo0sdPyTqmx0UTQN/0KG9tG3jPVhF/mA9AsPg2pJ7nh5Xb
QcD6epvwb1ED74WJYAbraD0uDKsrVdn9L7gglCEx1HF+9hdUkpHdJuYUa0woHlwY
08Fe+f0wGbLtUioCg0sm3aYnHWIh3DE8e43hxLM9sjPYpY6pu0PBNuk4+vkoPAAp
7gaI5IY+ELLPgYMHY/ePg17pCyTR1qxDyVE/DNhVXycQ9tjJ8QYS3jnpg8zlwWXe
wo5IyIkRCddjecgIZoqb5S3Noqn/SCE7CZIjM0zcSv7h2Nuz2vKeAte9KAPPhRv1
LJ5189+MeWpIyiIakENAwS51ckFxc66cRRa7Q2Uxi4IqSI4wGK4IlJ9nvWK7Icd4
bZjm32/Xv3OYczz8pn45CIlDV79IUYUTAUcXs9LXOytSz7fshfV7bWYqycC4EjdG
vOoaHBvT/J5wA2Oym90splJa7s+ZM9jVm/FbjEgqN014jS+ZrFLHdtVyQsA1y3pu
xdPmoghqd+oNZthCTXRvxLuM5HswIl/mZWD0AH5gww1vulRXgQFseaF/2TwyvpEH
9pBaFjRqMft+q6VzLvXyZw07IJF5ASmFRCzBDDmqiQvPqbYRo70MHGea4MDMN2QB
ozmTy9KEDaX6rF6PiArPy0gxe2Wnc0lm/5FjJdBEhWqeh2iCUfhUjHhQIPASICwG
FtFDEhXzYkRkw2T690oLICuNVi04SRDW5P0Gt3w28QLv8RWlQcnmHUL8Ln6cKccP
jD/2tE/5Z1cTt7gJlSEYXVHklygRIZMVYk7m6/70pBLhzNIoBeTlrw5RrP9szkU5
MvVgoM4aToOoFlhKS0RgLJbyjUY2YYFcMUwIyDftyg4trjxfGYa2Z+sCOcR4R//Y
9hEk1R6y6cvk7LkVcvrR9zVGToWphl8mWpFdJz8zxL9iEXZjSnf+3LEZbpc8GW8J
NeyevFmz8FAJ34LGnlw6HOxQ3uny4LPGRPDWPTs2HBHg8Y3Amva9rmNTkQdh5NOV
9EZ2vHP2SgHPE0oGcasiEppSANdAvvplzHGvT7ErNJDmG2VDqbUzzpkPQG/vYgdm
FlgfvsZGRMWUa5hx/eAk6qSjW7j+Z+MONyOZBE6/SIbKfX3OXREP8eSivUMokqrV
s8g2oS/phNLVIoIbc4DAygGcuo3WOWenxLatqzy5NQRNW9OFvhqxxo5spwruxlUR
ddIojyAsq0kekQkajWHM1HDLM+aE3IqefRxK5FxAE59Ggg1AYD1ck7G5j1xBzkPT
bZVzcNafqTYA6kEOyu8MadXw/nmiWXasrhJuv4HD/fdui/ee1zFLxnCN5dmeUUDl
HVkfbCljusDkXeYFcPszWZlNCC8MYN0RiVH5GqjTbiIMkKJxhUFh8df32n2S5OYL
DYSdXKFk2KYDq6oJsELCwHHRadxU/TRbRjfKkdJCGamev76sqB8d2NbNOxgBdGIZ
75bTetg4qtShWr7nnqnpL8gUTGCURgQLGXAjoBMwp73D4br2uzTbrXZrMIXEuqvv
EJpRPKJYmlyBPru525Aq4Fn4Oyx9tQANa86u9GQfdnVhFIChzoufVtJA+7DOhiIb
R4WC/10aUi01ET4Uc53AgSU+4sDD6eU9jLgYn1Eg7cUYYEF53qj9Ph4vgS+ezFTn
RL7c8qy//n7wxyh+UMEIvnG8Cg+6QMtxcDsipAwQDWliyuvcRZAGaFtmue2Oorrc
fL1t54z+ep+13Q9QxlsRR/Hqq3wlErx8tL2QpISs61lSs8HJKl9Y77ypshTQ1hEq
cKfXlTCNpd1U7M0OKDlYNa4+Y6m2okORGXIpcDv8K6EXTeVEYRvx1ezTCuBzKW5u
1LPXyE2ja0VehOeiK5oM+JdKXPQky0lzJzhlsBWUnkDW+xvpsvuN/D2TS44Xruei
N+t39rtD19tGaA3bL1Jfk/Iqslj2lvaDsOhpdE6GWDxh3zWU3rwcnFEN/CIUahv3
/nojyIRj1yBhmvMySLEqHyztAHBixpuUyuuswcO9z5NM1vRz1WX/1FaKr/tYtp2+
rh97/lFoiysPT+B5RAY4TpPkuf77wow1LnVmgqV5aqtq6fDy7uKyQu0871aaZa6b
Qgg7fL/EDCP2Ar1bSAw1SytI7+hlYUXJ/yQYZIIjDSOwAv/KKSmGiq94cTvEEf79
vIqPVT/3ZRyOohg7Wds2D6Qeu6bGEhm5yRxpnj8GMwGNFFQdGij5j+avcJVoRwsm
qm598es6r2Qv9pk+xIr2ji0xERYoqo44YelD8rX7ushKUEV3YbaN8uCLgwxy4jv6
rQtDVg//qsaLt8pkUy/IGS/foqXefaTzvCF9hPRmPTlYA49Dz74ChClNAK48SSJw
wpAvIakMerQ+kHsAK80nCQcGfXpXnRD+YRUPK2ETScFJXFHEBAW6k462OsRXbrWv
ieGAszYz5lEy4o54dsqd80/ea+IF6BJCOf1PiYlfUy9Aj4IHRp07Ujdh0MugRrVO
mdGKMnBntr5gNgxtFdXV7e7pg2/lHvlExLV/uWSJjif+FU6/KMpFWCuOSi/4YmjK
E2Y4u+bpn6X4hIG1BnKOrHqfQUczqG9BGwRQMQJjat/wdV6PAtKoriaKMu+ww2+h
SfWtas436FCwyUGfFHormtk+KsxaqtHRoxnoTb/Q9a6g8XC5FB9fXErG6RGurfOW
J82FJD2CpWN8sfJ429xif667/iJUxn0RoBHHfE0sG9R/avtwWA2YSGRZvaZAfgJV
pnLHRoY8tpt7zY0REi+scv2Tqz1EIM/AhOanHNzQZY6L86pX1Ng0fjSscmJdSIlv
kGyPyHuj6cnhAwJ5lpcZau+4G6OTkuv0RL2/HGhDVwsGfwBqhx6GiUnri4DdvuoV
QhYXAeCFHYYMVS145dTOcKhwOkA62eCSzdizGMc6YJBwqK3Vu+l8xX+2/2z8CWhk
2KM39cjhgrN/4lLSvDH9STn9ALENwIfJZAVj/6wsq8Y6YLOIwEIFshEOfOw8+LdG
uX4JbwnFncdpr35HvC2mMa/LT5RVUHJPAffrgtgEPGYb3aO5oQrvos89GiVAh1cZ
8Cd8Pc0xE4m6sVKJpj2H3Rpbygsi5IKdT+qXsJI3bS5EEOKX172vPx80sHgiKFYB
jt6bMb1/vEPnC8bvUcPgsweDA/UqBnA1YavIpZpMC3RWzmkEG9hPbv0Pp99Nr0fb
x4ZC0DXYbkAWouTdbdMhIhS5bEv5HiJmuNFyd9+P2yKKSBG4EfzkciZvDZQUH7GR
lkR8kjPyP4i4LklJ7vO2GFF+a8Wq9odPoKJQ0uInIpJlKwYxyVbu44YrZmSYBZ7N
uzceQIF7duvs69P9xdUFfpBVg3oPHfBH7t/g+a2R9iKd7pEVAYdN9NbuUA74LN9y
PxERkp3kQKcff+0Sv4Vml854Fv2myffpXW3zPfe6oL84WPs1FKIZhFFtWocKRGne
vVnG2tbitxkrjU4YByNrOe9AE2tLyi/ZKCFR+K3rel0cT2VA8kO18I7PHaiEophM
wC5SkQXcyQ59hZXacQoLkvpY9JEr8F6wq1TzGxIkf+pU4UUxTdU1pdlZxRdO46af
s5oQQ89xMF0c+O9cNmLTIYrL9alQzox8Wg4Ut8FL4ZzTJhM+G7VO1noJNoA64f3l
pCWkaCBlM4URiy9pgfzOaJhDOuIX9IT3Yf9APhIbKewInHIc84euNSnWKmuH47iZ
hTVigxZcq0QpkVEcYSFRFxfdLGIFYhY5FaAxrAw+tPAZrbyck4UcjWhBPdOzAars
7KKTbIoZ+qww7/aCOsvQXnvUOFZCcZIwgCoXnoFethhqrQS+ZGjD/ky2sRNftJYu
NLrY4fUHKCiVas1s7GgWjsE8ZlvHraoV/Ww6suGxzwY6DY0xQXadaTcIKSF6UeWw
l58fT8A3+I1vma98cCyVnMDDVetnLqLBGiv0UODOtLdnuWl/jRGrCUcXTKtLdKcG
53k96Vv/HafmKH9TqxvKOjpQ3y4XxurrJwVWliqJCeBIyHcDBt5Cco6MAfpBqzGp
v4824bap/KK0pZwiZNJwBetvAd5VzIXiPVF8EP8m6Hqv57a3be7IsvLk+NRw+HQm
TPeudz9y7I39CYSc5sDSJc3SifwCQwiBxA8eJYkpSutPzYj1vW93J4Dj3oD5xV2l
8IOb/swwAdV/+6b86qcsFvpUBi28XR8tfilpIVsmcRqaQHnFTb/LoBwX1X2g79Wa
IVCesqwUlqO/Nfh1b+22USquuCWEAhYrI2GNfsEoZ7Rbof2vbscN21yGy8vQTKCi
1ITvBl3q1auogfdjhEOCjyPXTd4BSD5zCuiROEboAkBVX/FctexqDOPnEU/xPJ4y
cOspzp14bhwmI2eoX35XfkGIBdNQkkALB2gmD1CnK0VopCk0/6DMIJRXMoAlGoRA
vV1d3zseapGMjPtAE12jeWHYxCwUeNVQDibhXhoZIi+5jIelhnJmU25lQLMqFCy+
MktTzqDCiOmSYscEmv2RgFWbA+I7ddK21/6T+hyHrGGpgns99SQY9gmXUkWZ7HY9
BidGhPfdTq/9Sd9o304jqbEw8ovaIeA0yOkym5RdkdqGgMw8Z8YBFFPUXkXz7tko
u3qEa1f2ioJPz2XkJIDYwne0816/RRkZm6mPjCp757lISKwzYofrCBMYcfQ6fvk1
ig9UqK9DngsjaCFxYNqIJbKTCxpK1ISgPDNN6MLtFD2hqRS94YLSCiPuYKxLJspj
OFlQgeVuNcgRQ1KTuGa/rJ9VqaVuuXq+zNigZrBiX3mbC1Gvr1XJ1v/sk9LEf7fs
vP/l95jRW6QcF6Bp0rMfnITJTlkyF2/8W5lVglu9gVKJIA72tlnlUTLGUUIjlsOB
6vf4LYe0rwSjVdMuU8OK52zlsjCMJ7iNr1l/zEkK8rgc5FQngwQeMZhhid8tUdXi
1eofm5GCSvN9ogZ8jeQ3qSAVETkYmO+chHdhiL2ji4ahKwnp5iA9GvupUYqyvIhG
36fpknCrv7q7FHCkYYKAE9Cl511hxvmCoTt3T8iLRiDmyhaJvn/xxcRFSqxisvC/
aQTZ5Tt7BuGAm8t2UYLGMCAgUik6BIcE/IvwdHi7QA9T5bU4XDl2gxWV8AKUiswU
kEa+kKqeOy5DaUpcSERzRl2QbK4mJ+OZHKJW/otrabC6za+MyZPCX321hRBMI1mL
p8BLBvbyxWO9j8SmoYwjpFP71zUQj8c7Werdr06jhxzMUKpqdgovWYrHmc0wxgNS
q6zqhNBYTSS/B/K4vcgl7b/0bu0NGhY/d5NGeBjYqqs2al+/ZM2MZWM3GJEDXnHx
JvWatDK2vf7rh5C8WCz9BbXW6qvhbqt41YuWp0rDB2EAmlY0Qb5r/4lbRKJCmq6V
kffgYrnPieZXFsiM2xXLgz5/jCAb4Rx4jwciMEFv8/NZy1H6AGJj8dwLK3e+h3ou
ODq1XApHlwWcq0XShcdbMlqE1SjzxBrcIh1MWgAlkF+Gd0YSAtHIS99eQLf01Hka
d/DI6bfsQqHlUgZfX/zc0H4xSyAmSHh45GE9HvbgQo4gt3sYozPTTsJz1E0djbxL
WSlTd5ZaivY1dFSyK8kWmWrj8dF3+DLEMcLg/KMnb0pbizKkDlE88K4dHqXylR6l
lZLVHjt26VcuNrsFED3tsXB4Yh7/x9LLT2Z4ujNkr1qAfnHSSq8sFzaA2K+NZDYF
o/m7BCQDE4fn7vgRdIqD8jjure80fCd659f44s0Ti0YFn5aRfUn4oUyDMvJBcgNh
v0Pk8hQu7ZgLnqS0q3vCx0KungaKZfEB7FD0UekfVnDk4Ubi6X+oamhYvaRgwC1y
tQQdj+ARrgt5MkWXhIQPL73j7kMPndhU0sSfO+l6lNdDwAVOXDcrfdWQp/kcCXvL
eykNil9SX/NOP2DynF4j7IbE8+ukJfFraEpduIOO40rg+Yh1nTxIuRm8NoCjxD97
QDQnJKq890NI6Ip4JmE/lboZW69Z1L6i1Ke2QQ0hKCil8RZ7vE6m2K4yCu2pqmkU
YY5ctPBX1cyydW1Od1M2f/damcVW31gUEGhHfEYE2VpmiVKWFvF5YVh2CPG8UoD1
pBf5TIpPhfmQmvgPmT7wnYjE3X5OcKUx5WmEZxl79BToDRFRBpdODOylCy5jf83f
XOQ/+RlB2VmMTb/hnU3asu1znhmRRWbLis3zJrxGM1F3vWGT0FPkAc68G9XrCRGs
KlrhB3McSJDhnNQcDXs/RdbRKy/QPXSXAAFfcxPNcJEZbofaJ48AnAN0kE5YYgkq
BqNOja2JADI14Ux+u2+4/uiMo9e446vgOj5Sq6GpRNQAFpNZNlPUzT0ei2ZLkep5
Qp4hrIuiOC6SkYMFLTIBkFIlk484HFin5/LJMIqX7DN68A2YQcL+1l56+HE2/N0h
qDHgFu5gokfvo2t2uSZs9eW6PktfcpO1xTcoaEyglL1wBAeOmrGvruybSVF2jKGw
tTPBuPYS/TRYyqfzMkzhqVddkc2tokdqs4yQUKAVjAZeFiCOC81bxyi0xR6vteKC
MXV7nkDJftv/zxK86qZv1LMYuqDQkSM6dUorOVk/lWO/Avh2syLgxxOqzuXdemMs
CH+4hVBszYMfNI966FqFq1dFq4wfWjzorG0kQ83sH8paYY9KId0A2vPDfDw5T83S
VGEiOVO72msg5zChk86RigWMY9+Z0j9tpNqQm78CiiUPA9JZs+5ywc1q+4Kol+1x
9PSF6eSEAMLiXf0OCwnaJTUkvwa5yvIcyFWUQS3eC0N8MIxsZC84Stc0wOP70LT6
n5dTL+01IOxd+Lhy6LxdAEQvb2TjQ8e5B62c+kXoi3yWR7hC5lBrPOu7sXzCpIgd
JXSqwVvGbN6T6L2yJ7zu/kxKH6oN8m/2AumYKHvkYuBK6FlycIBZNb3NSQqSuZEE
9dxvJTOGfJN/NTHO/bKZZIW5UT+kyxyOLEUrdd+GcFzEXqMOq575MGJ2Agn48qOy
k38b+UVNuLuZfP/ge/rWsSKkUuKZyu0iU/1Dxct1QXpRDGW8MkFgXhk5oQCX5uzF
c8UvbWuM7g1GIqFcLVQXSweNJIHWDENuLFblHWeG0qn2E6iKBxDtXt62DNRGNjlW
u+MiL23WjaIGzvGEuz+7nP8MLLUqd8OSjTRl+f6RRUuxt3JR12QgwYvtBeL7d14I
SfUcXAzlNNovtLRSenDlG8IF1Bs39RtObjj92aJSYejSqrw81QP4sXkLQNGTqvuU
vZz1VXLZqq62DI5wPnbd6bT8ZhmqqyeCP6qW0Vj734hO7l/BfR2OZ/kxJTKglzaG
uceoH8gAvZgW8OwsH30eFZ+iaKv208FyQ9EPLdJA3IzdaF7whxjoi6CZ3yZRhKPK
aOyaaVLRLsw0mas88jrVmAlsWXEDlL+na9UKoyZDkplHdZ1RE5nKRQ3+4txLNEOt
ZB+rWZnCRHFY9vsjPtO94gXrxbz9JIzFAkkqeCtoTvokvl8U+TLn9FeQRHN7b9pj
jcT0cgALzhRCLmUb627TVOfPSp90YPp0AXJnc2QoXQda82iutfhUJrogXPefeFlO
ROlwqpIYm3yK5M1BOduNQ/qp6iCcIP+9+vDd6tH195b7XdnCTedr5CU50h9xWP6B
DKGX5Fs3Wxi9ylTBaA32bEi1fwHlRrwcjtj74BtC9oNucIWYd78jHUZBV34VE8Mi
cwd4E80G008HV6mvnY/fE5UAm7rFrk5JfCo8V3qMYGL15BZuVPJjLcIHfqLD9Xk4
ouFd7v+Vr4Ki33i6qGSq4itSjUefSFbk4tvXWpuTPVoazvLsTKlJ9V398mhyufU+
aB0XEUxSYWmLX7ylpMkqOn4MTDEgZP/ojR8yud3rc9Id7n4sUbvfLZeAeFexLiZg
iww8TFHbBatAh0ix+dshUSwX4XiZp+65tN5Xw4gFY9rDYRnEIgx2Z0fq4CtAIQsz
RgxAAg4JeSO7bcD6Cu4LeL8nIWdte6opP5FOByHGMpwyVsvRRp5rqjn/NmYLXMKW
aBdNljyVSFsNYIcPEI4vmbj1M9fIXPWgwm8U9E42Q4MaNTuuVGT7HFbIcLXGIRv1
jd27Dwl2D2engPTnJh3ADoZQA6eqYElT0hHRemBWSrMsv9NSGmOkv2qVCA62Jllw
XUQnKdEgpwdESu5ehQfcUH2Dk62hJxWClDxptwhv4QfoOiEB67Cfhcyw6qwwJRom
FK3LOnwlMcnfEgLcJM4599lmH6825iyyttMHCY9upDcHL38WuxeKtPrbAYy7X52g
bIM4pJyhMCS/twRt+6l/UmDdz2/94ehlgPw7U/u7br8vUCBEF8eX+5G6K5RlZgsn
6RhKkbnjWPUQr7y3FSrFC7Hj6yDUvKtGFyv+F3Zzg3jj7VPfRqglrVSUb/ozRfUm
VfgOnnjqLqBeRRq4nUdzBC/OcAPeG/94kKBs02qGj/GwfNnj69BhgnYLwag5L496
2ys2EuzpHiDznVy+taKuBsNF93S8JJuTjQRl6iO53ms7Ytcpp59nNw0pIJxLzs4i
5U8up61Vx3C09hvqPAkD3PSJivLIQ3ghMDST4tQTyn/XN7FMI7xQT9AR3EgM3zW+
c8BEwATZ4kSVEy80Wc1kG1SkV7S4FhVuiP54mjf8HOYYhZAfMnBxd3Vqybhu7z+r
eVFMZ4W1MYgIooorKsOf4qjZ3itu7IWmz7s1lEn+843A24WQ+1I7NRoO1bIoEQgu
cA9fPSsFNHWnpVZvznxPfmUfYKzRcmC5y1WyV6VwBqoMLLYcuROrMnndYeyxKl6C
d/j3A0o7v17OMDdVE8KxrmjyoQ3uYfiyGlWe9vw1ShxQh8DKUFradmTHzzODRN/c
tjVvaUgRV5nuFYYFGMmb52mUvRGhK7z5WFpSMaPf0CP416GPNRFzLft0onMmgG/w
DNV7MCSL+Smj5TyYxehRe/87N8AwpB+2J4qD3p34B8ae27uKAQ6JToULidLqlg/8
C3XvxBbsClcjcb1SJG4dTMwSUNrymL8bYNG/x9EVoNWKj9xQHsIbi1xhrgmdGpMo
WSMwhu6LJZQpzij/Rs36Ks1WAKSr0lqQdzjymsXi3hFjQQb2wkoOvK+rZXA7I76Z
gOvyhZsw84S0rKygPUBm/J2/lhpBcoLIxfUunfvWzH7+jmjvOvZ5FI68wFDTaNl+
S21rj4NBRFS8UGJkpFUvif4XRRGBzJjiA04AOu6qcRJ7xcdw6R4iVkK4AIoj+iKv
Ty5dN5pJ1HYQ3K7G8N8za45Cmgd/Has2xxaBgyMnNuGG1h8voIxeLoygSZS5XH+X
C5BJpC1c9gDJJb0Fr1P69lFhIvLrlIjqorIi/6dzkbJPccXmnELuTiovaNVZTcr5
sxIuQK4LcMG9p+zr5JNksyObfxHxRLV4kmrgElCKxdI9CsrWYujSarYNZ7RnzI6V
xjOpD2hKZaLmCZJdgoGU7BW4N4oE/Hg7bvim+xEHOZyvl0nPgYuksGaaWUPAK124
Unh9P3SNgU8IqUF4YMrnpnh3u5kcvKLKbalZyrQmqCXa9cffxDuJhYHf8oDHsbWr
U2sgoXQQ42lh2pZ0VZVfP+CWozhSPSVIlxtHXiBwrTCFXRO3dCrPsaptrrI+woKE
wkTkjoW5rx6WjTa6kzzEsbZWYeD+sRmz5HK4d2NlMz13pOsZSSPdVLsxiXgoWqQn
a9LQ+FKO+pcr/jNuLL8F8cADdb7YKnQvgFL7kUzv1xLdeUtvtIfwOCj2iXPGEk8E
DLBUV+6rJ6EUQoUGJ2w9GkKXmeRfXwAbNdMTtTh1cPzMhOQyXYHt1Sl9KNdZVTF9
8RdFETWQOhNriOBA4voK6lHU+cbybgsFNa129ymwjGu6KY/Ll730q4fvXjDIvrms
fsXdOLn91J6rLeRJo74AHwB2echxI3zlnZggjVTQ9iw1/kn4p0FZmT56ZgnPntF1
NVOjrMsoBer6O1iMb1yUH0OY3K+VACgG4PE1KQPEBQJaQvZasLSmr8eEIAuSyxSf
JkB4GIg88qvz28b7HEPh9BnTffg7CHa1H8KiiqJWL3ZZxvKUwFzGNlMbtY6c2H72
6W0Tyo/AI4w4KE6t+89pEZSX60A1v72vwWz32BsaFktwWKcZSaFDGvFr4eN00yBv
8OV+xPEVfseJRIsROTuQ73x7Lo9djwuNZIxWGN/qD5TLZhtCqgxxN0baKqsS/TRS
4+c5gxub3M6RMHJtrv4kH5DLuEMc4G7WPTATD763vq1QsXpJtC+c7gMGNEfZI1QW
ch8G+uvNkPbOyX4pJUcfZ6XfpHWtp0Efkynzf90zopNVIb+5bmyx/P0kYrKzH9tH
4hM7DgqR6VSm1e3Uxkg8IgaPwN3XaajzqTPEb6P90sJZitO2y7hpxeFs5CDcQEW6
jTQsXmd0fx9oo5nZhQiqP7Lp0+995RqE61ygR2jmJb84RE8F7FGihgS70FbhogIw
opmJLn0yFyy8clV6L0i0iNUTpm+XGqZiZYWUdM2PN328Q3nK1sednnzt+3hHsr9K
BAPcFOE69dldsaPmMC+UJxiRM+flsS5tbSiWKSxUEbySyQ15VaonKGiwkpn1tJgU
hAj7WFuw33X2zOBlGPou0AmfRTVRxxi7FnAHQ7A0ucjtBTX9TmGzC45pOKB+irfS
XgvD3B47JZq3mtn8L5BPPs3R84Y+TOv3pEhQ/sSm3odnj1tc2UMvyDWIdNH0Bm3U
KgUI1E0DqekqPRZ0Y6ctO74zdxtZ63+spTkf0Cxy7zNS5YttbIfz3TBH8yzxGbOg
g6oAPhxmjyR4bohnXAKfJAM4y/a7j4N/EgFvvGSxbQfqcA0ETjWQwP89oU9Kwm9o
LZ9RwBVEnKjliHonTm1Y7CnZ2KkSUrryWJzdlER8nFWkpy2h0Vgd2bp9XpimMXjO
Y86eNKbUvjAfc+DJ3rf2gOj6zNLp5e32u1l3HJI3l90Ot890QUadYPTa3DN+iUeh
A7pAjQUMrdsEkisofj6+XZtx+N/sQ1OA5bPj0S/rH6sdsvnz3jhMixqYyx/dFHNp
BQ+ur/YVFFxQjxBtnxw0rxRK9cKyIy7b1NtHIXQ/1JSy9giSmPLXxM0pjLrt93Wh
rF+NCZiCWFYnDUJHHbsFI1fEMU3Boredvm541eZ/l2apyVvL8lonT8v/5sddUBI2
5HD1N2IIGrey3g2bX45L6Zys18wL3VlyZSvKpNdi3J/DJ/9mLlw/DYAhmWCsI1yu
KgtQlfDRHG/mpEZs3Px5BJo8xTAXyR21vfax1Yf4iWw3c5/nowsi0zKoF9ZooCdY
/MEG7zh0aZiNqZ3sPEk15WuO5JJbzNbAGhwtv8G8d3bFI+wU8qcxLcTiDVrtRruT
GJ0NNNOAHdGbhESBGtmzHYf/m+9W7t2j0OZWkiQWSjD3LUZ9RH42RJNgURn80SOj
i93j8+/ME2iaRwvUUpj7sYU/vJKVj36NL/ZV8ES+Wz4zo02R/pmgjQqQeczS+tGO
hpvujh2YJJ0ecKkSjxs+BCmVvwaUd563YOVhhAKyAsLJ+S3qt3zCDrDGOPyC/Efx
0G/T21ARE4pOX9AvkTHBec2J071IEfBCsCCgn3eoOJUMPkio9Te9/WRAcjXXhu9+
Ml9zyQXOmINVOhodDxJ38LYwa09NYQcHzDvtQw0/7OCtSEVTPbIe0OAIwUfnOf59
mabbcHHr8gyqrqNuHCUAqyxuDcrujCryk4bB8n/vIaOrZNZrrGwLIRhku0yPRYtu
T2p90WKJvlV9HxE2GneNyj2H537y2e8OELESyuB7Bmu3mJwZcr1c8j3qPjBb3nqe
cGETzB4zwP6sbpRHcEdxSEupOf29niOIGpowhT8zg4APzsvIH2RaGL2P9L9U2vwd
WA4q9wS5wYgLTCSJ77Bw/3HVVbNrkECnhsUHgwvXAXuPWdpQ9ZDDftWHxCABMxEg
xZXKG+5UwYRZOolPP4wNe+vWUtONV5jH1wxMOE7zsjb8vy6N801s/qE9P/1xrKL2
LAiuxdXtk9WCQqla+L6pp/ZW7tEI5/dtgjOzb6PMcdjX/BXwKfZhdnKnYt8dO42L
W9No+LXnwDH6q7j+UDX4keJI4SQ11zgamcsonq5Psdmou/B1AQNL5yBAhYbbHnxX
1cfcA5ajCNf6khkTBuyR1RfaTv9aVkJ9mA0rQNaq/q7hCxxyuHS2Pnfp+52qMAUf
qscXcvPywT8jiBK00ZK7fXKzzlzq2a/QfqY4zneF57mO8vfCP4txactXNPo5ACfM
zpqwhnExvbwCpyq6m5UjGztu8OBKfCGGu+jioe0KWMkljN3xOlC6ZKU8nDVM78Ku
0mY3sU2Pxv1pzMS8uF7GSsQ2l6AcK67+YINnnmrDD9I0YpPVLGKB1aIUe1RXL5JH
veZ4QVmSoU7px6LC3iLw3Ph3kG6J4gMgKmH+VLksY2vZADAtVSt1ERRYdBBbUrPZ
CbnsaZjv4h4LvWkXLc4x4avRZL8HEEsn9LYDxzyIyLfsm/9hk4r5jQv/E+UwVJFu
7cKC37pIw12dEhWvT+4mC55Jkb+a6Rpv8gIeV+SZY/vqNnzP+OEJ0U+UZV5DFURg
uB82orNo9tcs0RiP5tSOu5wQB1UuQaPYy5HvKWjDPmpUQNmh5iQ3tD9C+tQkgDqp
0bpzWBtTNr7mCGpN9oe7wUN/ctJxrP1fuIXk08nBQr7IoAsojDOUbUA8H6OGBe9r
rFF8HSfJXVehoa/mk9I2WFddDKAvSOW95PxFabKF2STjKsAVSh/jKPdhMzoMiGm0
pmJkwN88tv0KcvutU04Rsqkb2GZpskpTeFTXRqEN+y6X04lIxjFIe6RHl3AvJ/7u
33ykErwAfyaMV8C7VIrHUTyGxKFdU4Ss0Auz3Z/I5n8ESN2zTKxXLmHBE0vjOTkn
SEeal6+4Kqugs5Xq867gi6UG4a+FIypIg3+ahLewuq3jkEwTJ/zKlCxHECT58vmf
MaxmHOoEjArUSDilB0iVj+Tzy3rNTyBFuls4rmhzNkhOgViQFDj5LsokAniHnes6
s1dbe37kXqJjQdKeboqEzMpSKR0n/L1cVE+TEvzz0KnGQfzODBAmTqjQ3w61j8zK
tVaM16ggMpFki4OXPO28UBtlqlPCftGJlhjBJC2wiZNlKgch7iwe4KBZwpzMs2d9
ypzhpEbX/Jy26KUzKIh74OH0IjPGc2ZHrqjQYuU6LbkEQJ6rMgF1YzSjNXYX+/WG
7qCgGJC7BRMglmj0fJ1iCdb190hJZYusUxKTJNE6MgHMUm/4CzqbIVFaN3FJeBvb
/ckBza3p4p4MsGOwnxjRootDoB6gfZfMhSDfcbn7s1fKK3dL05hZjvL7gSZs0M/X
FNcf0vnKtDZNUiheuTQD78LK5qBunF8W/Ayw1Dx/PRe9yWAxCYyrXJl4gyzFE9IL
ru3OZN0GFrAdfsyA23xzDYxVhJHfUJgiqPVDNV6o/q7Q1He6lMELcnVTjv/YP4s4
CzVYo3LNArZO7KzonQ7H0PSNGgE+7kUw9klVLIm6zjjLQQ6CcRmPjQS/YnmAFdU1
xxMnxoYB2UiNUjJjnYp+0jXNycdOKmjQwImcPSExduoMR8YqxbW+Jubxvh8f+GGh
Nj+CTO5QYTsHSOGpShzTs7DXibLnbQdkR5Cf+YlYBkcTkJiZIjKPQAfHfu1DZy9y
cAr6dxzwInkAM2LtJI+b8/8woglt5W+P5cdoD4PUqdHB548rfneLeuee8GQkNTWa
MWjXhuRX1fqjQn3z5mbPlMIaosS09pn8sHqBpNP8QsDRpm+691+fc9Win4mxO+Fn
xyXVb7o82tN/7iU1Md9m8Y6PvjG4MI4uhT2aTemuWtb6mxo1jwkDpXLZiNLuKr5R
VV2lDCR3Sxpd8dEahOWFn5t3SqDpum8Vtmkhns0V0Pd2g8hOOmD3xh2M7njl6TpS
PyQxL6OXWYsYeBCtqS3CQLHDIW7n87wrXeR98G849l0cbVmZZh9E9HHKc+cj2+uz
JGzAWO61N4hJXCDVP4SRH1Fbc49CUS9+TzK3wHMuxbrb7LnfwjqDyFOZcss2mCs9
xzfUUlHpTk+Zj9IgLV2ZUZWjGYCx4DglqB1R9WvM700NbKkthoXQq+x9c1euWb+R
jSZPvbACSV7IMjzTAJ9cpF0vxepYVh0zqMgRAaoWRsyrh7LhC6eRG/rRudMkIRwW
+ggQOEMTxmsiQ+fIg5gtuVabZDtjDfvYdWsYDYvBE8EqParqGKvTpFmLOSb0/UDR
0W7M9odiy8qbEKDhKjWPyLqMIvCTQ8Hhoyb2WTlXtZmH7IFIfT3t7qOVpGqxj5GW
mEWlkteiaoipX6ksQHhef2jcPDS6Zc0wgZuSK/oXgGhYZvlJxGU1nx6uZ/HemgyQ
+9TCKSqJGH9PPTCcayZWPWcC6Kx3bFSrk6tUqojy+ice0vk5MCx5jYmR3lXK/dEp
J3rnCt4mZMGBwdXZt98vU2zW5DfuwdPHzOFKWzJECQGCsXsR5dUJZH+2sncZGQMp
zOl65KP8FA7z2HFfTQmAZfyXCRRB1nQ9jsEzKXundQSmMfnSK1fVt4r8A8S8eqnX
a7JfIzwbAxLfq9iwy0NoWPEkV51POrB9nGa7SA7+BCWJXxTqRi5hg7tHzCbxEenF
dApcdwWGQc3QFVQ+hh9iIhABPuDHzea36wsvrgiKa1+cInSchURCr/pBSCI7Yqel
7h0VHtX29KnypSmj+8eeIn6y2YVaj7RrTY6gaFuPcPMu0yHGNlYUrkvhE19LHEEV
RIR4coaqi352VDWiKKHK3oyAkR82teB+ifoKQesbj6Q+4Ofc2Yc7XLnBY+KKqo08
Xu1saXlEgZYu4n2ZbE6CK/b54A+SkJutf2KXJ5fcgcvcM7JYkRo6N3YSecV7nKLa
PHJKgTKGCAD67pQIO9qkS66opS11MBEpSYLRpGSOLQ+vZ4Qfp/72wPIh4GhCBlxo
2plgglF11q9I5mGYAOvA1GgOxUYmwFJGR4LaraA6DJGMovAbgjyEV2K1iuo9Ewxm
vTBnE7dXrBhCmmGR88ztkTf1W9TKPznDDrHz00RJ/nsuWW4+HqlnT1P1842f+JfP
bYTSf7D/dWCu/eqnbvYksfz0aAPDUW3JLdru/AmRbu6W4pxRcTNIDxF4ilyx2pK0
wPU1t2l14tLgAPa5ieDkFM08CwrSA9MJi8qr7UdBmkrlkQVLk6zbmbeM+TId9tcv
+rn/gGxEX8dWq25GAJctoGRej9NEALZYQoeTjvnxLf4YY4LNg7HlCJG6Ug4Q/VBZ
QkZVbpepJIP3fzgswDBqjndw62mjvUB1hLlz3YEtmuhvKMTHN72KexRogJSW0OuB
ckJs5R5YW5UTyMTeWUIoMSz/5OXL6rG/J/AOKY1VK6WxkGaWx6eo3XOn2Y0H2Iz5
4zFOa4cyGCQUnjaOXLoreHWbO7zGDNcUFRojxtnhKLH9hXKBp499L+ZfwZP4ylXO
Jfv8VfZzELBzl3sLLFyYPnlb7Vy+G48pksDuND417OP7LDeCXHOKrRX8e/iXZyds
CuAJwFREHcehlM6E2yf6d9utD6ORQo07gxCEjHUbilQh6YiOo8t3IWOiWY9FBp3M
LmtYxOHmsAb4eDxHDBJwjNagqf9Ob7mpOLPQiBAMLE//n4H+KgGrmx1ji99FyX3L
eyjo9qgF8XDEDJaI3N5Fs+f3IPawD2Cmn769/oQpgiwNpngUSv1kRPp+ODgownlc
tu0TySPntbqbAZ3rNwio7CB952j8gamiYH5jy+d97d6HFp0Vs/JMWHDTBTer2ss4
/913fsVFyUNwJtnyEH1/EMr7UXALaL2EvKfSPE4QVidavjmUOt7rPHWSlxrUMZ3Y
8E2nUf4QZmsgUGTkIY1MfgFS3CYNx+OfgQpgzVV4EGWIkv0n/X6GOK3UYuyEZ9Fo
mfCi4y1xyKLaiGfHeWIMrektk84d+m4dm+axU+HlmlxqguvoBqDyYWN7duJ+SZGs
ImptXSjaIL0pEIZ/vTnDjAIdI3dHYvcWITSHiwmhclkzXZ4U+G7+zPAiHc2UkYbz
PsifOqU/LrzaaKcL77X4Ty7Hwl5s+7b6YKRGV0ubhjWf5rm0VLorbY8CpzmX1TU1
LHSzGQuYC0zayZWfNgAulXOQxNnSRge0DWn7Jv78v67Ap84wwumh8oUpZ+XcQBOL
u5/Gt/VNO2yoluz09P7GDDIrc+Lqhhi6MR/0nWCuY6wLfx8Fez1s6IoUITNQCja8
0g8OLKygTcXIbicuYJhj2gukmEfk++1+Yj1B6KAPBPAYQzIBfnWe8gWE8p3dHkdN
XoLe+YMan8pKLT0UJc0Lfspan/CmrqI8D0iVMMvCrAbUwpHmlmKhCh5D3Leoz6Ys
bOOe436rTxDPZ9SrSok2D3L6xaO8wbAiQCvQSPXpUpT86IeddvbwCdVvA02MevmB
xxSP7IvufVHVa/e+gECb4MAQaMB5JfFiMFC+wO5qiihMwYMLnpMkQpcBrdUFIXna
d5AJ8960npeqSbjVEau7v4/qNd0puKz4Wq6hrba7WiJxdD0QGj0S2OlUbhG/9+Sq
YJZVcAF1SbDqKW2mujZFSVjIDMCQfBoLAEfcAmyYWNrQQJt7fInjuR2+mOCS1tmf
GPjmmJyhnAJvUa3a5nq6Z+G+C5OtuCiqfwpMrFNiuyV6vsqGbyuR+2C7a5yKlE1l
8aBvxdQu/OVD9yDKSd3rRXnflIKjS+mbDUjVPf1dc8OVtpY1vyhjvwxI4BG6GxW1
nQyK4k6PPcSkcWxa+scY+iMMuBmhdQiNJGZccgg5OARHHgdCrzoRF/IF/uxq+C9v
qlzJrfXLRWcvG60rql8IEbgWP/1leblqpMxjWilUD8PR2PgzyU1Ri5ktTn6RPnmH
HvjQYoM6f46nzzRvjejwrcmAx4M9nBhu3wcnfUMmp7lq4EcEjqr2QuHmgAe8/CvE
TNDpulCPWyFN741+siP+ZYWK7/CwEDAX3s/JcRFMUrQ/jlMmRL2kvDG/VVeFEkxv
X7mGXZFc1dLBRj8Mqz4hn41z6H1lQgjeWKTGNPCd1JJJS9Gh9kGWg30kuZhxG/9o
XxKUpdkX71tymw0huuJplmjqnviyQ+sHOG9hYQvXrTtwrevHKD9TaGldC6U0gbhr
50/klvqUiW9LlljGHIeSTdOm/OLe9uQRJEXYF0Uq4dpObFC5nIdP9eb2P/9KkVml
ibcM+moWaZHb2jFlm33F75rVZOwkgGe1zbHbclmrv3YNYVUB4eDOFuJc1ubmkPuy
FX11eoNQPcB18efACImSiZc3vT1yXRA2UHh3obKQ4LJOHA8yz80qCppsK1hKiAAh
d3oxnZpvcgPdjJE3nqGHi4yBA8JqjYMPPMpcJnuJFE8czftiMHSbMaSObDaPgpCQ
3glx/vc9JFeDDgrkIwuD/ViRweqIQEUuCJgVpe6yusng3lmRenmKT7Ycy2H/vJJo
TIoIRbtzFaUT5pFNAgVMA3BBnK4P7Hicx2n5DZfKnxtII0KlEaG5/myzUjaoO5bE
UZfmiKgN3bDdRW5TPOQ6UUSEiGIHp9ql6iI63USYRx7mjLPdEMtBZcMviOH6Zq3n
bhldCSaKyMNcKp12SR9IgPlte4X2jd3sad5T7sUjivZ1EV+yW2Fbo2aMmajID42F
CzkeN6CJfve2hdPJjN5p8y5mpTRTCJe7aS7++vavPjqSC2VVufLHpmIfVNmT/TDw
linsog88F971yZchAY12F6G65YwSyVv4oN+L8D706DWi6sCVaBYK8fKY2seDp8Zo
loNrmcuKx+hfcWE7geNXGd7e0POwz5kvrPNm8e5Yz5W5D1Y89UkSYCCZCpKcM5RL
JkeInCI3kU8oK46C/yx6n3sK+DhqQ6v1DVM2nTyLGmKg1jR734XfEPg7PCWKNf0V
hAJFpviV9MH3ljPSHeay1A0t/W1+CTwYlB2j9yKSVLrBJ+1d+wu3tBd7lfnczAA1
pn+2RK8m4W7TcO7Ypq9gkOwIytwuAK454fIuBQeWhphGp1L4SXGHiMKdd/0tOBWC
cYOVMLsIiCmpaevuCv917i7DyzW1rNF7aWM/kXl9XLwCpcJ/gKLmDIAQ8ki0Lyel
Ua5UJiTO96HgU2sr34uOSG8yv72zHHo+EMSAjlO26CW7HpUOKn/2Xm5phW87H7+5
7ol7d+jQIemPartl9DGZRdIR/YRd7z0TnnZbRzwOWUWD0+nOdcLu7IyaxpOSPToo
PJ/0OLJCycYXFGgia1t6m32kmv0lnsJfDCGnTOUX/GV6fO+wFSuxLD7yKcG1X6j9
PvahHj6d2NdTWQUcR4P0GRrU5RpitS1LghZP90cVnGkea7uFnfVYkdfm8wQQttnh
B+q2+L0ZKO4UHASZ4ZvzUlcJVR7D5EweG2HMNC4Blmeide+fusyPFb8ScVYktMdb
NnBS+3iieSuRvDqM6NPXTWS5BC09wlZ9pMbH3chMLRWDNmHi9u2RY94T8O0fgRM6
RMYjFNsN/LWpjcg1GL96MnwTvtoNWFlUmHLyVlDw4JiDEoox/sVYcoHTTZOxHz6I
3tyAREKe4lVB3XwUWXRbUuoIdmv7kaz0l+GaBAzL8v+DMAtHgXMLkTmwMEnbgBFc
DtE+K3pCHExMMLimZ3Od6bfGZX8JIr6RWhpJUo4QCsl9cKlksAE4w/k/MkOjGa9A
/CTMuOLhPhx8b+IOsAZpRsiRpFeGweK+ZYYw3T2B22ajdkYrJWkAWkjSMHVW2Nuk
McmQ6G/3kETYIt3iqvB1/plpcK6nQTD7Z8uaAD9+nL5y2Zw+6w6E/BHVKamLbGnj
CD8KImQZ6pUxhdmhV1bK6fmV9CN7trmC+8ULhdwti9Zebk9mgK1AYqUGGl42jo2r
nWcOWSbMmM6MFfU+yS0rqemiAi0iuGr6Ko9vt+pZ4mRBwu+vfygELgko0r/nBLGd
YAY2760KFDVntc3Gv50rz7x1O+lLJMuREvG9obMQIloGY21lUzc3lWAxdptN5jlK
AzCPz79lWmTwW9yYDLIU945v52bcmu9T6H/ykMGNhNQpB6KwYx57oOLYgFkodI02
aZ56G8B9N8CHRb8kNe0hhwexP/PtBgFGCno93Q2vO1B4SFPPym8DmZOz2PklcDlL
/+NpTFsnuEhv1dQXlOsEv0hnGPiNkdzeerFuYas+6S0hVw7tzK8j/eLiyLaMZokz
opk8FNEpsA+wu1dBc+ckn1Zx0efz3C8b9sN6d/Sqcm3ypRegR54xwYTv1ekz7AXT
zx4/PX3uqgDScyddM22n7OP3R5DRHm92UAs+sPFR/WO76mnNGc3ev+V7JfSRqIsG
g+1hjGwTlQnU/6f8jtha21cZYcr2eYdRESxURTVgpc56rJ5iQHgnoCWquMWF8NqP
ZH1sgVUIcYFrepZpfFIkxwyQQJ2QCZIpJcsnEEYQpK9/o5I15Mu3Ksd7+gfvozxO
7ByI3mmH06HbtwdGzb+YvjBBu0Wlu9A/IlRZyZN9xmrt8chbYg5s7fJEIcqpH4xr
dHU7s758pFs71/rX8FsHdU7UdLNPBVeaw4AQdiHkIaqcrHtZD8YMPbRrhwA0GHFc
5OcJpKsmciBvvnKAvxR3ZKpFahPAquGmbRRE0Wkrdfb6hUrAUTxRm/uMqq8ZH2ek
YSrwt5qcOWrnc29xmCLkfVCO26OX42Svf5H6BjYjCAsz/W8BYhsDWnJjwlDux3UZ
WAcrwZkbG3NjLppWmA64EFryHBSQS8sq2Ls4T7mD2T4IKwvnL9V4USDTy0i+401/
LzoKhjPWoU4Be0Y/wDt+8mKevHHaEhdpW4RcB3UK886H/0z+HbTQaHyLenTokyEq
W4b4tlJUAHl9gd+DEnBYF0OMzmSc8/a0paRxfPT/tybRGViBbreCLTMKmuAI+HsB
/gzWNp0j65fONYJW3jccDHgFA9KIqet7/UkrfmppxRlyVt0n47W0/xWRVJjqmWug
e7Pb4EJ0+kC7SlVVz7U8TRUgDk/IMb6rFfrW8i0Yvu7PKMfmi9SAeDE5FpKIRnaf
gTVxka39gMSl0p5X/+ynD7F3wpDyNCv5KRobsxhAJ/5XQszOAbpnL4iLY0n3AdvH
mroXzgP9pWSO0oS/jJO3DLNyOpG47uvZxPgjXUY7WzlE1m+9tejgqTTSH1fWD63i
rdrcywhCiXplgyCZ7tJkuILW1YXsKi6HBbRYi9i4hwndgoU8syQh9vpeZ9ZyjGfX
GfBu30M+xBLcU4M+7Fx3q71vO+V0ik5NpbQgU4/xiOH+c1bjFQfoSLHux9Cyvnfk
9Sft9t0u6EuqqbURd139HZfgMox7B97ZYQgtHwkDVBWW9EpWXdR9DlgxJ5jKcpz8
zu036ZmUOujkJ/8WL0g4CSzELKV3RzyrkXnMZ11XwJ1E1LlSTsLe9FB3cT3iAXUR
Wuzou6jKGlhQ4EOfWvhCy38zZ3eJEqrDisz3X1U3p9edapwSnWOfyaFQOigf8SQ0
9592hUgKjgn1GWgrZ1YcSwqN03MCLNMHtm4huDJSJW13ydhBbNLvjHOot1Dxtrv1
0MntuxvL9SRCKFkitLzajpRH2m6BbF/4KaGOfnnwkGhjRXdQMUkmkFwZw2iJv5UI
zVSjKts/9zDqTVJPhHk2YiH0w8uZ7LOLjZBXg8n9tmfVI2i7XZVU2CenfVrTvo4J
sSH8cwWLtFuYZXFk8wYoyMtHDqaDu8CYrasU4n41UCsyY+Q5EUjh6iEURQfSvhBC
TfCtD0LOdd3nl6wKqgjbg4h0SUIeG9DH9VupNTIzZnDmqF3rjXZ+9Yv5qLchV3wc
Z51IdbQqneJtXJ+6IwDYKtd5Fr9aS0IV7lhXroEQ8Z3N7t9ES+MnUPSiVMc/R6/s
5Q2p0+PLwYqAQ+y91gcnIroKDxwRDSxGBlhxhEL8ewA+wIVd9ry+obOy9/D/IiR+
CrMSMWPYo5QInPTOHU7192cd/w7FnNv0MDjA6vmmydz7lQVJvmqnwHIBJSjk0Kns
IKFT/NO8BMHh33k6R5QzkTcv7cwXj4/M+E1PaD0MAt4tnwAyYrmUbP8TYouB2nnL
SubDletc4+OYBKQ73AWAdBg0ORWck9Ua9Ottx+AIxKk8iKC6Npv5ZxCqFqOrUmBx
yOmynQNEmsX2zjpe9Xl4VvEfLJcWclly2BCBFokJYlITkn0AO/myhkguFX8fJiry
bvI3x38ZhqZ45BXg/k/IOFCHLfvEvyOQb36ut4vy5SW22eJ2KDutBzUCkcHArdI7
2wosBZfKo8LycWwao3vBH3gUKtU8qmKt1XL6wDFto/kgJXxb80NLQUd/eVF/M406
CT1gstdwkpw9I7L4p0qblgnl+loSGuv3pm/IJaih7m0CqgjGTCwsEB8ajmCiU0WL
3R3GZy6pOITeDcSDLH7Pc2gCew4faW6M95DwUaYsOIU6xGPHpg6HWSZ26QqrN5tx
muesq+xCZ5DSnxPCe8LkfHD+XoqVEbPe87f2pWrT80BdR8P90TZn2CJ8qRD+05LR
RQlijoWWSDQ+ZjqPzhIxtjOWUsp48dTKlKS7M23j639kRVb6qtdDCGnfrLPuQzYG
MX9BDkFdTHWMWd+WI0g5NGsShP3E8ZsaibTgef4ClDo02nwbAAREoJhl7rZYlqWj
d+WppB03GIwd1XClQUrfTrSbqABHTW6H6ZfUZF3twqh2U7ZegMrRY8+6hkLQGa9u
89O3ftIr2OUGOdpuYiurfC+ctSVoCKD4JNh6x9T4Ku66ryC/q51Q+3WEjEu5VqUh
A8P3zPJsmQGRcl42CvtMSg0T4/Ljq1Bc/4pssG4Px6l+FWJtnMCC9tsUeSkfLxyh
KVQZWBNZtRBOOgzVLz3eJQZ67nlsGSAvdv35p0fCBszHSi24k6jLyhTWU8aFOLk5
EH0pMzMmKqnpWchPblngoy/Yb26uAbzw1XhfXbWsNKGSrpRyd+xOIC5cIfMiSLsc
P0L4Zn6XdqrGNxlsXy+F4y6FxfIdeOWWEYpTgUPsWbF44pe753WHLCPxbIlAmAkU
HM5Zg2o7ncahT68ODdPEYAD1lEpX+U5NDI5Oal2nAqvkNsjPbchmii4JtY8jaqYM
gZOwz/Xyk4EvX8MIg6lPF4e+fVaKlrujKyJqZW8Jie6rEHdxwbQ0JKYzR7YNDU18
uBnLiuCWYngBFV6LaRmIaVPL4yOjKW+6gRo5BXiTO6XV2lmmmm/pDSSOPo5tQXPf
eTTLE7I4dBzu1K9eINvooNAaV8nS2JkyvCg0EAFMxVRITfcqk0FXEaH43nooBT9y
5ftuJ3GyU1WiepOdrkzu9AZ2are2oDRLK7oZ+BxA+k7XexHAJYPUmGnJ75sdKtzk
7/Q0T40rWh9VhY1Gmx554VXfDbjQepc/R12fZ1PXAogbDHbBhzqzzan1sRifQJV3
iHLM69I/esEA9iJy0MuMczpf4+h82fRGhT77hj26TMtpXrsKOVimUoPgd+97sOn6
Bk96cPkAo2L9rzRrO/Bc2VUsJd/CXB8Rs76TZJIUBngkbwu7L8Wyf74QSBxcWe4x
c+FriUU/cctaIs1697mbqUxva7Y239XHM5ow/He1KlWPUBoGMbHwM0s0k8Pr0L34
oxCQIui7zRUGTwgz5XlV/Px+BmRQtjG51l8Nva8ACMJZZnkym+u3IsnA7L/AmCoR
aweBox29wQk/hmqnRVwqi1GVKTsZ/bQydKneM/diExqRlohp89no94t7c3mQmSP/
sIxRrLE/LOgM4BFYl6dWQs6wOS68NtciHZ6hNhvUhJM7/5XBuiqBF383QHqssKek
XTX21dIWirHyVCyGl7nqbkZEWwNcgYqBtr+7ktyujB3LekvV/CPb0TAkV3V1ubP5
k26blL/yt6WSeFrrLHsQ3Af4VILcVpZkIMIjV+xx7ZMpn565QCDclS7eA23kSGU0
9o8K5L2ne5EL4RKxJUlHOJFWl8aI+kErV/psYllPmDv6Y7HIAFBMWAGPplgVGFEM
JWnkQnjrn7H8jeZp6A4KUpV/qhOPDIbsh4X2MlPJVqncyDIsQSPm2FbnNd69e7Cn
RKjSaRVCae7s2l0oyLBbFnJ64URp9XoInGZ/8gb1oHv3bcurL7QDcjwUbJqXZyJ1
iP3d2ucupksNQUEhBWY66KzZ8m3Aif2bCykB/By3kl+LutfxgyxM20h8PNBiYXhu
wDhJquywaI7Tn7/5LCs9w7HD74fcyEioUUZkr14hlWIkZR7UsCpNrNfJcDEwjPFH
Qc+XH9HU+vwkZ8txJRrELfgI9INexjoOgl1oS3xiZuFp6Qcz5oRsI/yiEH5tQxYz
4ULvBEaYydUL79GDyb1Wm8EHqSd3itji8Z6qHwIkJkXfomGNcxOvzYCYQ6s+XUIr
I1r+dLBaDOihsvbyRaBIguDu+z7sr6M5Fj8U645xm5cRaIC7ug/7wmc21GdwCfRn
A4LQvdQruu45yANDBlfY+I6QFlSe459SQ2iWYiZvV3aOzpA61Sr/9IL17bUPlXJc
AETLA/Mv4LL2Il9kL1pH6f2aD4+Etyz9dORfUgOHtBq4wiT7IYnG0vSvxRIiF0iW
vaH2m5MU1NEwus8BlEPQFar18K+2vDhPiiaSPRJdx197hxwV6ntSyzeInTSo4EC0
urbj+CARudEdoWRVfGGra2ZEjSP+lQUiaRRjFgrl4c0DxTdjXWbJO3IK5v9+rLFh
2M1KXdkmafstEaHOiYIej17JdZqJd3v1lyslunA2yBEXud9I0bgE8GuloJbCbUvp
41MqNzbw7Pg+raS8ZpFCa3CqkVfnNqWa8Ezmw6iON0BeXpFmz+Uq4yKcw/tnBpBt
2nPGk9NUXvsvqYEFGUnM9nSXPtCRo9VKPMRc29mr9H20CBwqBBeijdhwlFSCOS3F
hErVW6RBGzamLO12xmkXGR6+zcWL6GoXk7wf1GPJYXeJd20TQePDmzQgFonGLF0f
hTOQzbrAY9NdjQ0M5DDtEwHEwNscHfAaa2lJgzWj4TAF7x8RJlMXS7z4MY0uUF8l
7kwsY4cnP2BqLZmQFka02jYD7U9z2IWU47FIE2V22cR32x/YKT/N6A9qcOcWlsbf
aj8zUuFY4tLHhWDbFt8xfCs58XSsowVQU1v0S15AaziTYXODsWbBSH4tDowO9198
LUcQiONJOLYihqGCrqLrkENyJFxryOI5BrtBB7ZtelLxrkNFBP8vk2qVm/9rcVgO
0gXYwpyd/UYmx69ZColdvc3PBZus6qwjPFz2ehIU5S9VleujoPGhccN4JEy8586R
xw3Qs/tySthhw+ZxKZYfcHLTCvJeyyZFwjfl2E+hqXvUCIqN4M1VCioIh6xeiDza
BZyqJp7nHb62uQhhG3KC7kh4SqswqAfcnRRG44DAGXnj1uAW8qyHscBtZAABLpbE
W8jsxwaDEh/6VO7wOupvtUV6HzDmAi+CUP78Nh+FJvZW6BbGV+k55KyIx5PoHJ3W
ffHpBcmLQSluVLjNRs+h96txTmK8SOHGP0n8tcu6pBFFoBg2TLcADroizbeSBM0/
oOGt144JnlKUFpgyG7IehL3rkLPpknFfLze3T3hZcV1BlcqITz2i5R+jUut1Evvc
x2SvwvlDCzxkDu7D3HdBHFO5eEehGq5YrCqDAaqlDgLSQxoyxPAIyf92rOnzA2vo
8VX60fIMwJNgvv6R5dcChuAUvC0jhb98Fi3br+8hJ+2mpVwPJ9l+Bph3p9FdcLdJ
Z3Mkq8MHwz1KQmhWon3qGCcajJozZGhyvHgAFvNPkOpqp6lHtXAKEcP9D3tKzHZd
Wrlb1MUrWH+d3hSEvFyJQTp8xH2WhR0nME1TVNh3vNIYX68dLbRMgsbPRjhvvAU8
CE/TtcWe0nDVmi/RuJWUB2MJz4uxQ3Bi4+L/T29nqEYovbSfM4r17WRGteS84gMo
2/zh2hzdPNVYm6UlYssU63GrvPrcBb13uvejwkGCEMC0E0g6DEmLCEojIt589ILn
Y+hkqeJTesYHRHv1sgUT+NMTQATdfRCHygXqE1QPZ+oTuAOVwF0EnkFBm61WSUHp
W8lMqpS8TX/AgLe7ZR2806owW3HfzWjVeVMwP10tprR24s6vynOEcjKqmRy6YMey
HMCoAOk5FuuRq5jigDkkqnESs+D4GvcVvNBClZ3Nl9oZaNl7j4i+rnGFFQXbmvxo
/Fncxq05GjjGjHEqll/5fdjMFdAxmTcI1n7XK8u+2qDJ9DgorSRSULIbpSvvSOuT
ymryzSl2xHUQ3skXs+mx1DGoJsd5aMDPX/EhttkwViRHXzB9/pHaJdpgX+o44xVX
kqSQmaGQkDtUcBrzFVEP9U8ubwzyRORw8I9skGMiQOMUKbn5mzNXJVY4v5hmTvj0
IbMQwoN/qJ0j7W3m6BSV8llfT9PbNSVv5klJyO3ZY44qKg241UeEnykfF03mhVdu
9YnXMailzo+uAt8J4hW7UTnbirR0D3RsNUoVn+pyDB2O2358QHn+ympyKtmuPO1u
RtuNJ7sDFbiAtdxuiX7vLoV0KrpBMa0/bTHP6KRoBTSIJfux+fjHAiDQoZo+qMjh
lySTaIMfzGkj/rX1lPOOlwqAvaFwnbCL1vMBWDKQEM0ym383MSIq2RJ9mQFgPGgw
KL57Jxshjt3sZ80r2vtY32p0wn/PfrQruxRu8l1adx6MDCW8R1665ADSuGBRxA5Q
2hPaWxTGueZ/aQIf+wm7PK5xgTCjxx8OQBq4ZtRS8kwzJ9W/iGOhxUhYxvP0tn33
8MBiQ6UigxFvuZ72W+sa07VLyzDIz1zmH9wm7RNJ5I6/O9YiEbuo+qBdh7iehY2T
Knbe9VHFTKQPRs+6mEIO8VkCOZyA8Gi6q0U3482MuGuLeOqfAm3YIuGrO//+kK/P
QCp9UuYKDqONz+IwJq0T81jHd/rKWAP+UaBvPFtL8KrcKVTr9SH1OT7+bb+fBwYP
/FZR0UZuxOwFV/xlwyVRoU7GQA0F5gWFsjenkvu/gQJ+XGxlZnyTbiw3ZBSgQSjT
/E4Y/3yjl5PcDHzY0F/11laGTaj+33PKVdbdnMs6h3G69yJEhHLTJI7jpd92iUpC
GqoMnMd+diHcAmelEBEk62FtRikXhpd336k50XS2Mvlq1hncmyStyLkNMqapN04S
Ywdu3dLIwNMmDpDID6UD6o3ZR14sS18O2J5gymLnWq9ZujRp2cle2FH6HTPIxd95
IYVOFq7CRy+ULBchwZPXGUDP022BIofTSMjiA1aB6+V6XKFvkSflXbBIFIKtgwJf
FDNtUqVRuBjZohWwUu1AV5DVj6EgZdHRmpVLjjNUIyhMG+kBjChUFC9cURnRCp92
eoOAgwT6hUPAMVXkO4+6MU0c8/UyhmRxeX+h6MzRuCgBjoDnI8fLXImIrCXMGASt
JVbSquGvug6flmuomwvOnaRPzE8fI6a9ADlHPW3YJoO4ZMfpuNjLQzbyx9slx8vD
T7v3RIcUF8PdDtX0nciI3MecZvr494T9c+C2PW/AsT24jCWi5v4MAnzk96P7aztT
gSVfvYn8OxqkpiiB/oCzq3v/TL20wLYBqBu44FQMYcs7+I1iAGIH5BFH6qcUfrUm
magGEjHlt21xRsz8Tf9tCiLWinV3WoFbkrfHeDtDGmsXqDX8fU2SK8MTs366vacq
9CnrJ8SNJnHGdqUOWeC1g+YzbfggJtkYLF5mP2jb41Ng0bL3mo0x24AFHzylUv5F
COrigUoW+yFCb/HjDGH9Ul4Icn2zOzFYZUhYfyySLaXC6Cyf/qv8rkYkYF8moxf0
1WPREjTM1glZQtQoyiNPuQsfoTfVs/1OMar1kX3QeVZwfZ6AO95PAhlFXdMzW5GK
8T58owg8lMZgWTu4XfCRE2AhHYzZ3eSNi71vXwOrElJAWkQpkgcEECQ+wcxD62zu
BzP08TFDs5af8CYzmh6lzkNPAoztsojHZfJoSswCdUtCUegddNXeyFUBUH+8Qzl0
JQHYPSEdJvdqy/vivydNBE0V/F7yukvKhvGb8E8hunznXVObm36PXIjySzNPHAvq
xpSgbhq3e/e5v6ZQPD7BzrnUaS1vKdrzA053lvhg7LNNm9Tirg9p1jSHc8N3Vjzt
oDfyVNYTGfEfmr4YhhNfqx3ZMOs1Rf1UnKjS9s4U3jGM4UG/CcAwXz5pXre45Xu6
7PYR5LLcCui+Izvah6NPIGHitqYusImF6NBCK6ieXJMtLDSd+X+al8QqiE6k70Fk
M6MLrEqUSMPyoMA3R36P0/eizWNjlzGaOpkaOenohU/Fszi+qb0H2UiZAKFhjg7/
MveSAkiEgxEnqJx/XhHO4HIQH4io0W9zv9Tt2gRMdto0wgk4Yx6gz1AX0eT5s57q
bRFUj5auKndBz5G0Ci/LBc9i+t18JA+qX0nvCZigiUp00sjxlQAKzIBaokUwdD/x
wVQS7aJ0QxaHJgnQ4zkAS/T+t+x1iTy8MZ1WVSPYiBbMtSL0WaXfRmW55RUw0UsB
D7QOBxj7jA++JZgor6iBbCBy+fKB2YtozwzE+Xz09gCERngSCSP2474I7+HnbLP8
zVfd8/FQPCFNBEFI4bz5gJrkyCVaF8i8m4FKFhjsPsJH42rEcwOriJCv/rMrQ0rc
UW/UMnDle8hZ2C2d/G6NnH9noPbuveJv/3yLXvCVxo1JxkJnvaub2OFGw7Ykj1xY
BkUuY5IjWXirnDJTRQzUKTPBq15T2nHJiWl6ls8s4SrHTnExrVHVgC/aSQfwMRYw
3iQIHkxO4ZqNJge9KSvJSDVDvth2xgmyixf9m8gTPVAGNYxE6iK+HNkBDEo/98yf
Hlw4ZHmPMnczvIWEPYinoI6P/CySlk2l1ga6Ie9x730oNYSr3lRN7pdI3aBfm7Ru
1eCnKSgY2/ZfaWhxRkHHMrCV4ws0rEzPFm4klJm9KDEJ2H6l05V78E4GkZ3TsArQ
UgsTn67SExC+vHRs9mKWXA0wq4YSEHOBi5gYcuXrC/oYJEiWHMlw8ViJWlOqdFjj
72bHgJVxjaKWgzVFmUHLAStNt+i5hw1mIILM67Wyfk7CzJWBZ/RxhyxewSwWYdGK
fjdXl4E+vH8h79dK7qGzUTKgbcn4uPLYagNpzDkVo+m5K99ASIjgNchiTrP3iGQi
TZUYyYAfswpIizblk7Nk74pIno+WDRinwr4bKLtnSlUwCUUsboDfB5QdUgQChzVp
DqE8pSMzgVLo/ASC9LovVsfTOx4BIDqF63tkf1cTLthh6h2lWbyyNSj5eDHdbXzA
dcvPNzK0fehBA/zstn230i60QVO/OShNQYFf+IhRZZXYgO74Jat9cgGuCz1bT+B/
1axUF6x7Cs/3qi9tLmmXhCBzmMsuUlSQ2RmbUmzh5QpP/KVJ9cW2qC1NntH2NA0C
/PyYk8BQl70H8aXsKVrXGCNB0QdaJJg9Zw4m3tw1x+s4budQtTUhumi99uZFO8h4
onGGMqDv+L5HgF0h9qr0MQ9MhD118H/Lr5/TsRGXGUFMqk2MuujT57dle+LbEalJ
1VNsIPs8nijVWVe263UlfDUdpbynSOs05wYcXEVTIDyKcd8SzI6o548qC9BTGndo
PKdnLnsw/o9kHD0Ln8qxblDrf7R5VM8NCdN+haPpAbLRCQq4EkVCsVz2J+DWBWFS
yu24+K0eXBlZ3Bqw8Q8GSUup1UEhIpfXfXDeepj+wbfKLzK5MErGk15qIeL/znR1
JdAylcGMvJ3ymcU/ZQGWZ7/CkHn46HdQl+5Hwe5YesjOywchUuiMOPLNDFQBfQYK
sYULtvy3CxlmrN8I0+gHBvZzoxuCzKix2YlP3zaIYrDusP6HuUYJboDXKALEK02W
028qLj+bB0dmOEMS0f+8HBW4PCokBcN4wIPGnuNbnZjPiZLZTa24uEbZQteKLMid
j0VKkwHMP32kKg9/fBI2TgN3Mws9/u3qPT0W4dyZmCBZe7OK2I/4fyezhyCKLlN/
V2t/sFzdoN+X7yjC/Jbpl6ZraDZNuorIHYwxXKv7nhP7e/AC8r/yq+gnBDZ9BnsZ
rZXDM+u+M5WlQh5iGxzoExB/FCbxBPvG+5gf8OPVMIXBcrnql7qJJv+K3Z5i11E5
ih9JGeiyfthVkdIAukFz0lnzLU0PYQti+fM+sgQu7a+ryNO+L0d75bKpcuLhSOA0
eQ3B5Us63D81wQ5ed+T1pWHOdfVO5cpnLiyBFzxjxIqcJjkqMkOaSHVJmT7n4txZ
lnoaAipS/ug/EG6WawnaSjl7ddLw9cQ8CopMGaYPqvY+XdERbt9jmReQWSyLovs2
aolZ43IempZQduPXF1RMwJHqbwwHWoKgP6br8384K9v3+o2qF2ptRhve1QLK5uMU
CjTZVjhzlMg7PsJkKTtI0bmldm9Zqm1V4m8j7ARwg6LIXTwxjbkhpbBRjE7++5X9
iZMQNlBhbW6fK6WBmSN5U5qd5BmUBCfVI7hctd54ciDodsO+f+pPFpPSRTIVG7RR
e4kO7MY3wZ2cFHm2M1SWvXaNas74F+euSOrctX3lyHEshnKNm8di7qcZF8Xgvs+k
rYhgH8hInTZfhRhmyv3YN2SzfcfY1iwm+GldgVuOm9cvnCfRL2ynNN3+feGKezZe
j6PsIZ1QXK2hvSI0QHQ9D5yvIAxydnaBRW7NnEIWYSYvpHuH0NyYFmgXXZomyvvw
Kp4DtP9Nnw6OF+HUCXVHpK0vnTjgxBvPg158xiYwWq6Mn1nAPuaB6t0na+ih20hA
POwYF1rZcjwdO/buOqTXLdH5LpVA3xuNowXBJQFy5k7H8n1Q96y2YhKh+Pno+Eb0
vNGlBbqu35CWrdb6gQp2GkA8cf9XCjy5yJu7JMSX4kG0UhMZL2LyGzRO+VJxxBPg
56okKjporPda9yqOUeXaRnkTKCyFGks382U4opei5OINhTYPqn1r+mw5N8I9JJF9
xZEOQpIfYHB140d8lQXhwkM12rkJnlLzR/vRNpHCxJ6HTfsHpIpGD560/yVhif3J
5UtajLHE0v11Q5pqVCOL6peLDiXNeIKvauhdncWPWneGo1LBR21tSMOFEMXE5n9a
G8WSQRS0ufOAP1QqJ9j3dgEvip/+McG5iMt1pEdFXJiwgFFOUwKbPB3AtTuLj2q3
XH9zdeRcogajg8niWpa7hvfTV7vrJl6hJlBfPH0lgunvg7cgJ/3HyQHMmJ4gRV1p
UqM+uGNh08WluEblcgwo174zLLWEp2DQlbup4wbkCYaoob2iwUZ5ru+PVx3x2Q9P
qzDLyG8J6z2YVx/KlXzbiY5ywHoRaS1HXCKt/fRB5aO95wNJvT+MLVnDlT3odOJj
+j7UYnrlQLCmtEXQ35jtw5Ux0GSTVvmn6VCXwC2HEF9idYwrm2Vm2+/AsxHjmHZ0
QXFr5DxdvNUQkEFQRtmVqv/RRCU0k620ZmxSuFC7rTzgy2+xK+NLcOks87pQut3i
RGwppkujqGYgeKw6VV/Awsze0pzfTCj9kbDTDkP/GQnCToNf5a9YZUxa3CaDwPy0
k7Xit29vD7j7VYZwYS6VcocIqI1Q6PxCWl5oBLOqfw4XTayeou910xlgc8EArx4G
3FRvRdnFC2uGP2xpYdyUqZZ391AEPgfsMptltWQW3NxgJWmpTOafYims5cqXGBHv
2Yaqm6by4xNq4pEolfwkKQyL1YlaV1CcgcjfUFGXmf5pcFTWnFKuLIIpe66R+r8f
PhRg8btKulEqPXc1B01osiAu+dCrXV7rOzgYGqWWM8GT5JkNZRBJ7+P+mhjOVCmH
4wkxr8Cwc3ZUIuAW1jATRSK7QbTrqfrTVMZicg5KHaX5xCCJVIqGwR1Sm0bDmP2P
uSTMhcsPdG2EJILpk9p7FA7etZwWWIDbksixu5n6PEydiSS65Er++ib8IUTLVFG8
tP8dAouSrdQDAh/3pblDNv9g9Cl6XumwfPB22EP9t4/bLJjJ/BDovefBNeKj2IIW
6f3cG5xKexiCkNb9DGoKf8kvkKGmpMgXTdY76YybZvdgYIF/UuL8280ML1TckMb8
I6Dunn0ICyzH9pzAYEePVGedWvKBjo8LOygm/JuBkBbJa9NEnwqS8tMArcuf0W6+
Qm98dKVeBPKDl8RNNRqyYY/7uuk5N1L1pHrDUGnjStePt3YdraADoNU5OOZYiBAC
HrLLJNI0kRb2p+Ezym46oJGIuV39Ui0OBRia8WxGKm+L4+mCcis+3Q9pPG2RUxQ7
Jj5+m8ac9k5ZvZQCpbexdfFp4MaPD+dJpbeg2el9jzxF4IeibkVxShmn48l3RnY8
7kA4Rl0OApynLNkllWmOxhF6Vbc8Fhk1LPktA7Hi9WV/BKktvrtMAerTmvtLUGBb
2D+c3SMywjSNlR56AY5HiT3GUAQGM4J/2d5eOJF87qpvn+gz/Uz1ICbcjJQ9XNY0
vCqlFtmboosXJoYSYzgt/B1J2eXNJ8Yf569ZibMKHQXGc+UMK5tNgK4waY5WZOiS
CqxMeVMM6MhU0rAf9JJFylM4DoGE3YCiYG6plfIkBBefhzzFGqiVvPlWvWcJwCqh
7eMFfZ6SV5Ama04fyEO+d3dMFS64fJoTa861IRedpPsWnnjK/6+NC5WzXLI1h6lC
3Ir6Nb2eUS5cHOF9FqlG0FpjNBXCqhfx7LtpWkfJtQyEaNM4/kIwyAu2DbfQ1uC0
Cm7pkvrXQEpn29pYdlpotkjQPte6wX+a4QZnA4fAUoQt8b7KNuXfZShyC0GITSEB
LgTGq54xyL6As4S7K2hMucr7MTzVXJPTQhCRn8GLVn4NW/lQtndiJu0RPmD9alZo
ynYoy6AewkWVjbFTSsl/E+qWqkgbNIz0ZAQ93BpQeQcSdXmf9KdWAQoo2A+sjvCB
Sa9Yi00soTv3ZQSg8BuNKEfURfDLY+4LGGUD1hUkfGevR32bf4spDOHQe0DM5FPK
OPzHAWALpDOs0p10IbZr9m5vQg3x+4nW8c4V3zFN0+mhDSwxeUrfs18dwsjOxzrn
phpvk0WIIAffWkT/u5uX7Hu23bMUCgkOOg1rrVcT6pyutZXCoDHbe6sMVQEDhlBx
on0cfbkgZwfQZiTfjLudS9MAHgzBEDMKQ+16jT3L+igsVX4nwFS4tS5BICoPeDzB
qe3oUW4J/fDI9ocAs0cpm+oezuFmDcJmY0tLSCnJPI8JEqFCv9a7FfPzrVy086LQ
gC3xE1qCOQVGKApcwDTKfYhrP00+TgfiGUN8v6VGmzIn+r2NNtOl5ESc6q2ql+T6
Q+m8uGYXpxx0joldIltCZDHoNuU+IHEVVJykCmX9bgozxatg1cq5SfAf6MajnqY6
ObTSmffeLdPTNeas9Q9EaspqMJT15hqcyJ8E7rUpLx+HQulMOCY6S5NUCqHqXpju
71rwnZL/bRZFovPd85tLAi6zHCiqL6ukgM1A8EP5mq0bRHYBnC3yHsyLvQ543pNN
Q52JnZECZQMyK1HP/cl+ShI+h9MeTN+J/Ob82aGwW1yrt85LuVygljA/M2ohHJn1
iZkQaJOs97iU7WTItKDrrYgrlWuoEeUOPFP70EPoxx1utGZEmiBo/9NsrfKS+k5O
LtK8SO/0IjPYigDwXrZN5tvRu+d8pu6fJoCIBgiutup9J2wQfesctdvnmwXkvtki
m7syIYKgEzanJiT94ze5lV7E80SYfj+4Uo8Cc90ayg0HT/b+q2ug/ap5rN+qrT5W
RLxcKxiYdTfw5u3nYBFqHSzj0j0Gk7AoJTuVBhdwB4bOzLJHjo/bu43TZ+g/09Be
gc4QVH6E66fuIHmWpO8BUCnQAYe9EGYbfRZxNKpGiwVJZuRXy4Wdblcg0up9CVlu
uNnSm6uUmpkAQsDNhsoCHVwUsMsfnjOS4cYSPXgPxHqFA9IMwVef9bQCN3C35xI2
/aAxTjjuDDe8NcLfq61nFET/LvI5CX+siIKsKPYBB4TjrhA+qrRLLHVlNyW5jkHA
MklpQJBQND1XgUIyftP4gJbHpv59QWnJl2b2tetz3xWhStBEhcT9bnMeqVDTmICP
DGRkl32btgatQUcRc3fZeDaNwmWMg+j2hIvbp/Xjxbg6+uyvHN/qlEhn8l5vRC2Q
kiONqnCfMTJ5Zvx10dFIRSZZ0mHQrQXisgYtH3FoFKApR0XZ8kH05JUr+4P7uQVV
WQ+E8vZlKkCYooa/GjnocZKPKq7LlMOnf2tXi3ji0znosEpq0NQjPNmDYVb3B5Go
7NY1ArHJ1Ju2AeDMhv7VrsX1rcwQwZTkhWWXmFoPc0UeaVhdNrTKJA0/B1QzDRvp
jOdOSsJdptRER/GpHOdCxGXJXYGKy2V1HLJ9OSEbS3QBe6eH+7UNUqNKgFAmeRHZ
X5h/WZeL0ug42N5zyMOPilbQg6yn/MEOVhtSzMqP8NRGn+FgmLdCdxaUiehjHVt9
EaPNLbYnNCibcVICiHGFwyJDzwb0QJ14WPCLUxSQUC9MGaIGi/rxmypDtAyl4fRw
DBE5Qr9IwNq1CxPWZvKZjYI3Lc/jztTBoUuZluPvXFeMKEdgIFbbykJjnd4UmuXq
bWSw2eGCQZ2sIa7rukONzjY+rOPsS2GWbz8kPCRHnK4Z6U2P3UplJZJguVfr2M2p
0+NGQyX1FwkKHZbYQo12B44QU208T0+vgQuazuE2elwq/eKRaUmaBpxVofx6PkOO
AuGw6dJjOKHdTpkH1xBVdneO7wqWKe4BD0l5m5RODQJmbuXhB4gHvhorX1PhPiPY
9k0PmUUylk6mQ4+EzrCSgIiZ+fT+FTplQUOX2m27JdBFRJ7+QAky5s/7OFIh3Pei
LfHOEnXYsG93iM5jlokoxq1qRs2eGc8JGoocTLCredbgpEwervAFrX7UVRZom/1h
VmM/Yy0E83yokcNOJwrTkwEpbBM7z5Ql3OY57raH/a2iwitHRDON04YEjB33Qxcf
kuoQTCDJ30Ui/dUVe/ylMWgsiPrnvcmnzWFJe5vRe+iHkaPM8RqU1eRfbXB2D9/J
6v83Oq9/dxRXxnA4tQ4H+q7BhniGJ0bmAFgrdbhkEFcdZIIM92C15e44kE5Pwmcw
vS78DnJCMUVt7RKfMXjZ/H5CX4A9b67Mwy6gwJPw/Si81D6JWlVZOzS47cIuVHoJ
o8SNTDgKfR61fmbASLrb013oceWygmVgmlRmqpkDhPNvsfBNnJNcrUhGoydDBRLv
+/aJrNuZbqpMcGQ2Jxl2cdzbJbC629GTqw3k/v4iPalhkl3TFVav3C8I1eU45xt6
zmxLhdd3giTvRzkoP3eDmQuMVVjVL6nij/1copetiYrnNgsVSFSjhyfv6yRMnV9O
awz5jKKk0y9wwiKZWUxnlS0VoP6iHAvTAeGdP4JTS33f1XguSevCRbyw2NuZ/r9L
y3CIqMgdmy8oKabQ6hFG0HEKpNQVFtWxHO2ON2nhTiJQNhkLGUS5jR9uQnb9Zyc2
xoQaQHekpyaPYBuV89NDOCIPpe8U4PtxLkhSZgKBN9NdtcEZhnh/HN5UwMLgDuOj
9Ro1YIBo6b3LIqSEbLjr/cGsSMJJAdq9kC46RwAv9jJTHrt4Onk3U6aEHQoY4h/c
rZtAU7GWTA6T7byWYVxcN8j1ioHMsJZUZ9gwv8baNWrVnanmGE1ab1nwGUHK5GU3
nyx0T7vacpSMsEK8b/xS4hcmKijR2febLzY/laFnmZ4Kgn9UjkhH0nU5jmdjgJP6
eyG5eo8/RrexZTaasQvbGT7urL7V6jfYbo8eZdgoDTNDyaAe0x/BSrmuXeWsWA7c
3sJUdo4fkHhvfDWpsFAzrHcq99BXlU2jlbnySMa+OHudMAE2AmFi/jsSTBsKYZ8b
+UBDKU/KIGrsGko+Lunpd2Vrcn6HNMAwsZFQnGDOATo5xq9uA9dZfV4blAzkjhZe
hurz6iPmFpLXPYbNDDx5ssOlf8U2XoeL2sDpWkkpRY8dUiuXIUar5v3RN2ReYSF4
0f8ChKDbOStW/WdsRYgYkjOqJiw64fgqXgSvuv/hDnfnISHU6fTTA+AogtOf7Eeb
07Eipuy8m/vmdWL2SZh/fxyXrOLpWMvV97UChWwCrcwmiyJ7T6rHEqVsz7+5NuLO
pFR34uylawgll+FaCDUqPAi9Dd29FlMPcVNrRlT64dY8hh3tyCZGRTV2oefaxCyF
K5T0QW3Wdj/cs4UlRUBeXJ8M5mYTmchLuR2yKH7QSd2+abBudpSxVdRvB24HKKvc
AhgRNljrKsKzNk891QFthptGsVjUQTu6nZaKfbMK2DPZ495XmBpo19YU6uCguIik
O2CVsfnGZadSkvyH8QZ/ZVwU9V3qx+lj+pv+xHSgCgE3dxWPMRgSMfME2XijXDfm
HVG8h/Z1NhT6ARF5zo420ZeQTeygvu+itl1u8LXRS00W0Zc3IHkLCah5QivXqPX/
p1jDsvyBo3mSx3S0+yAf/bHFhvLewvoEMovdZyHYr7v/EvlfbyUNjK43uEEj2zEN
seHh/Dksm1mkLB0KlQhgb7FSNk/2gss2MHaLvUn74TrEc1m1zYjvBciN/JybsF5m
32CnG1wsr3SQ6mYfxB7A1glQzdro80EIBzaZc+2CbOLv2SBx5IbR1T+EZ/tNQMjF
w3y/3+nXUUub7wJa6jIukEKWNCl+LV4dbZuJYAqi1ded8nqR9yShKLJ6nxhZ+dvn
+sTFvUdJVMi3HCHOPmZGiVYWrAbS+aS6F075A4Se7YMHa6wwVTFuio/BlvJGncuq
SG/d1vaiYzHMykppvvo1MWuWp+lKmf34JKGwKicKmMwioMefmNzfY138zo7WoXo+
79Vh4oO9/7lJEUC0W0eVKnC/KLYYB8ScMsn3LfwDB9xYyFoIgf4a5XPlQ/d8U/20
YZP3TY4vd2UDUWqG4xwKs14/PPN4dfzkYvZjFaKsqQQqhkJzozfZLtHAT5y6kJFx
fle1ul/6BdcKyYVuJKhfZe59VVBYkZ5BZMR2+R3uDsx4exbBgX2muzPEg62MNxBo
QDeIrduJcJMHorCLVkwRyUYCWuHVOCn9dx4kS3p4DnckTHrdOUgcx8tzBvFaPgGB
PEqzUti07CF8NRtExQsj7I6MzTDUdEpqxynGAKRlLV5GS352oET6CsLGEEzkgmNj
aIne8ih51ZjO/kpEPDkyIhQk7SzLoLHIUJuFDRFbau4PNQOTZ6wEzACAF8oO2Bbo
8FZf4tH8EIl9bWG+3Mze3f6E3OA8NGrV5gI9oC225yGfrIxhdxr1kUBQyEDOaXOf
obhKo5b9Egcy+f8tAr2iyfK1QJH+ZpxTkA86femC6sM3y1MokVOrxsfhW9pCkmEu
IUfdUTWHEZ+kTNJwMT4xS3x/QdgABxF95//fcAMsHVeLD42MlOS1aRM5gJmQRla3
4hsDau6GVZJ+ewMB1RHwvEMqL+iNZ2cBj3F/AwIx2NDz/yDSAbMl9jOnyu/rPJc6
yUxjuKYidmZ0F502kEqHT79NcJ9oDZjRpgS5Z82nBrURoXXQ11Jv5GGbAzyGI9Hc
TlyLMGyYwkGyqX6X6pA6MtY/ms2xjRD9rVEA73ZD6sJdxeyEaKfepFa48PDqpMko
wosAphpWNYBoxVRQA/Nu1EWT2bZMFtTRZOAqCSpMvdjBULZHgo6gAQqrTdXHubsO
WAXATgtZyXmEahg0PYCsiC7DTUzJUMYSRWUwAIenf61OP9kffFoCG+oRCLNN1TmQ
runiIwtnA3DnDDX6BonYEvXYjh7XWB1WFBuQZv4jDixbpDTKFhaeMbG7NXrES534
9AuwOEzs3nMFNWSWv68gbPvx7TRKadZOg0H4DFGlt97dKcgw3gbGlpvAItIeaE0Z
CVhPYsM+AUbh5edoivNOWIp0t2AcQIqdwMBLpDx/zLnws/Dz8jK05yl6sSac98PA
ureu5Wj8Z8L5GHOsCFE5NXg6WA28/APs2Nlis533De0kNmJJ6pebFzY0QuwHkTr0
PEpZXkmDXE4P9lsBN1z4uxii7AJA048nWoFVmpRlfMFmFBu9FAQKGBrsBBXByRdc
nZxYKXYjD6cWMOtQWgbPHLMdxTpj2Ckc2poWrpcEKNvtJ/NlHo67ySEhQ5W8WLKn
PkDsFeI38xztjQA8sod8pK5hHOe3n1+5oz1DsKfa8UvVDU2NxbcgwekZ8yd5NRVp
dImGMm/j+dOaYAcVbVpcJvyY/Ptc9h175W29xWEtV7JH2mUTwdzFZ7GmlHSU4af6
UDXfhhCwUgbY3BoCp7yqYvf9S/HK8uA8uMlpt2nyumz6yZpvpgoyGVtWpgGb4jWV
5dV0l9fcktavp+j+VdJYdlTwAH6pYe+XOLzQHEjcxfrrox7ypIK0o+KtgolzKyh+
4Q6zi1PhQvhvKfGcBkDqTMeuMBh2AZZGOtfe1ssEEbYVXSwMFL0bSOb0kPJQURmT
7mMiGuh8Tlhb5PSISL+gaCS2gd0Lm/d1W3y7RtHbadbnvXV7NX4YTSw4crkQ8bxB
VZGyB1Hhi0zfH9bsTbuGAJ+nJ/xeBAFjm20fQmfgenZbqmoZZEaEXl0bxsEsItgh
O3MBoBw2vlvfhmaO7IvNZhdrqE+XiGjuIjAuykNJhYZkR2MUouy+YKW/hjWL679Z
gBW6vl8w5MX08xx5/YtCbggW5si7NFkHEhieEUrtIASg3OOL41Oi3UdrsE2b2A3w
pMbn2oJSAWu5Pq2PFXnb5VRj9jkt1wwPwK9r1QNZCd5hRgzhbjedseDTwfalR6dy
oaZAQlAnNqdllVQ3Z98n9YNyo1JZjBsZw+Uy0O9muHJD85S6AqHDDOM9lY8LIu6+
sJgUHiU/g/a5cDflpetlduV+h2YmJIr3FS8CwgRGa/jD+/+eU3CsUZRs0ttsypYx
pYVFpnS+4bkB+4TX9w4R3s3qkO/m6D7Ery82QyrQD5bbAgLqanC/EMQOPTXt6VBQ
FmF/5QoPbOmK0/VqM6i2rQmAWJBDCCRYY6Yvo/6cm+uVHWhHX6gxH3/NEh5jKSSj
MpyUhJXbLi60luPMPytYbMye7STpSitM2QfamXGLT/jbxiNYNUrwouRUUjSnf7Rf
Q23cQ86gnzHn5hIw8kVrKXzz4U9yMtepA92E5cb1Z+zhBRR7m49KVYoEAkne5OQg
j+7Ult/xC01YMTyii+2mN50NQgcYe8wnm47r4vYWbnbwChQXaCSHwcrOVs7+Tpss
1SgsPFaokTBR9j3zj3ZSEFZvSBAomr+ugtoYkNNPIvLPSDERwQhla95zpb3YTo1j
m4raK2j9VCgPH1IbGFQ8LpIT8r+KhNXGpdbahXww5vIKDEzTn2Yslac4G3ZdcmR/
yCV4d5kPkkqcq+EGqMfpPlVLCvrrBoxK1XYgYhrT0+4tPXoU1FiGY2vtW456gEMn
hArN/GYGx3/fLQhyldzHT4cw6msvsYx8gSJAI0zFAPsZBBJlYa/TWqwlqdGhukWY
5k81uotl3/vACQnIpTHfFbICgw/bHls2G0IjOJ6/oq/pRUa1jylnTlT1d9V9XmL5
ThNOznGSxeH6q86hbZOJTiymcymkKNJ4e+KG+DTLO8QpHd/8d54urvA5q7JCTzGn
kaGlzeEnnpuuGgYn6y5cqJbwzxGo25DwHhnyu+9/tudOzJsaKHq3d5GUgN1A90kW
VkO5tDgvXvq9XfsFbPV+6cxTMaA7Cn4A02tfA/0bHl5pQkmZPClCdWAojC8FVpz9
CAYQzBkKonwIaBLlhm0PCkhSK9M45iL7kc/nIpnVwnFz/qvta/QFT2wpg4xt1iwR
uCXhKLwLnkfMD/h92UMvCURzsWNl5F62B5u+ovJtdI3HgHYmCQplpFPTRpgTcJwp
U3FSoITStMpMj+dzCxZR9iPc6+Wc4DYS4jXNigtw4Nxvs2xfoTDRk62o/NrNugA6
XGgCZMH1HTcGtFZQyi6zRQkfEP2X5N9CaTleaB1Z4Cq0i6UNcJSXreAtUBXsRH2u
GmzCFknBLLYU1UmnorDhOep2oqyy0Zr1ejhKs/lUKUSHOxtGjtPQA5AeFJ+LbGl9
5EPAhUyIi6Ez+sNDiWdtuGnsHtF78BzLBDSJPQFFbC7LceKXfDzgrVBwDsQM8u37
iMPOIAE1y7857fFus0BT3/XwLsnjxjiAOTS8ext+E6ITV6xAGfLHCv3JJ0J9VpAp
nuzjRaxLjXc4zHdE+gDfWmQ+i5uA75w6nl0Oah81adt9+ls0Lm8alz7pbothK0OQ
6FKkZEUl+Qyo2vtQjSVSJLweq7H4Ut39yVcJelRBF0GXPGDDHLew+tPB2GSqFKXZ
5EWZcrs7R2j/iZDLaybTosg94DBHCdK10Oz09MXCznzAtIQYeyD4RiD93JWmMtuO
xeDuihnwlWWA0tbqiM97FoHZ1wG5UgYqUnWRI1LxusADT8g2dNGUp6lu1prrixQZ
gS8ZlBwCL3/euCAIMrEljdVXUHxCYBsvsR03yIcvcFk5ZKAQRp93kjO4YNxssPbT
ThBMI3c44u5bAvb/ZDp5rO9cjaq2tmGna8Ck3D97eBhU2u/MDP7LtahNBWR+I1pg
HnLrYJYEFMcAc44emxvtLL8I9Qy4I8s9VhZU8SeWjHJjfL/UqcoviOVzFEWO/opr
aLtSNH+o3FtbJrIw2WMQnl8WJV48mHlzFgULyhIPNymKmF3b+3PkfbJDYTPues6U
RxaF9YUwK6cKHCkw95gb0Cohtb2dRFJZeQuep5lrvK9MNnZZ39Fn5bjTSaouxVap
GcbjaGJ8xZF5YK1NXTrRGkF1XYpQ37myeuRJhxMhs6rzNyAMO4TcxgKWxD4gmbxk
xpzNAR7dP+Q6NSr3F3OdjsN0t7rDcpjxv4FurdiiClmBKQEd2Run9Z/POhHffhHu
jmpsfVP1Tth5IzWWtVxbvWe8jV4/DtqO+O3gETtdezQ6OoNsp/QVLxuN8kgKKIq+
6s8WiYWWczFPFY1AVwNMxcpn3t5y4Sn6AemNbqphR2SBBQzRtbAo3FZOfWSBCvJX
Ig9a/+ViANxayyWibBFN2o0w0i7M7ausL5ZpFGDO+z+Ydxl+1V0aoi/yWCNKFihL
tCIc/78wh/D5OEc97MyNOtQQTDZqlmyB8y3ZX35fRjxAsjjMIh127CqXrw7rtHnn
c9IPuC7vX9J4HNwYm3kR3a0AjmyIbhbHcMxMp3nOyXMZJnuztqHvn24f+b+Uk82s
uVB96UZS3C38B7jB36VqPI8D8m9UqZGn95hFIK0aQ3JMnP2W6B7YPZ/PNrIPv/1A
rDW7YEK26H5Rsl5eKdXN68sUyliqXJw2N4eZ2lYr01SaxxUgZw1mI/SJ1VpuaBHB
z3aEOh/cPQKczddR8AluzW3F4FjmdFfTAiI2cB8CbltSCGS1SxZj0G8WGPjIV6rm
8hNeSLqqa1VX4xUsOtFMAQk5x4wMhPhHs+LCm13EXGlpEalpGTxvMrfcgiWkUedo
kGX1JdKLPvhNNoBtcIlrpahBmvaXmwnq/8PgkhHtmb7Skj7Yxn6xH9AfBM+ahRqz
VFlpu1ewuI9gFpDBunnb4im0MSQJkKx3VNgf/xfm5rbkcbEKFe7aWmMJNjUasF53
kCdKFw5OW5rmXZ1rQ0oJynHaa8x1KI+ljdy3r/7hC0hT348ctC6lep/7wk39hjyi
RALdHhdDJV9A5TyY37okVcMy7/R88L4NG+QZp4Ig8k+GQbae9ptTq0tyOLkOk+mq
SKH162j8dRlxAx5HeRpNFoqpJnNO7oaucX1nRLajb1j1d/+tipg4wGpPHCWM3AL6
/KOkQcHoD6yPQWu7yB9jRV/DCVEymaZdYNUFrkR8XGWd5Om1bQkwxjCiOfORf8zJ
1JXrspQn31j5mxqFNxBBCAlosxX6Nd5tSeaSiw5EuLovMRAk8cV/AN2Xsz2h6+Of
BN14Edp8Y3QmlqssEQYcrzUz+x+jtTPYlxmqyfKPG8isK/AtkKy+beUneIAN9+He
1nW9lU/AtjJYv1WtK8DJr3dAyqNmGwJFOPVVyvbqUMFkOTfYlMu3Ztf+J1C2pG++
b7Oh3hofouBiRjUUPZdevJKwCytxJQD6ojAGCXYa8igfsyGbLdFhS547aSEto1u2
StWkzmjKn39BgSTzDjRWR2ewuCitHXv4pojAeAO7EJ2+pkTLCajx9dvTLwL7HAze
xrzlZ1kWT10Oe3FKFEGQ8b9GLJ49U27nf6aJvahwUaNNgxI5jfaHAu+tFKE/+Tkk
5D0HzTeqDnMUNTNkl4JhJIUkKiG4wzc/QfNW+U/ENNIPdTxieBz5u/F5Hpp2KZeQ
zWAu3j/Ku/gm49LRdSHcrOMRaXTCKlprA/BPIwXOMu+i1SgBcYj1/4+6AuMBkKs9
MNo0/63ohnT8F90cuGbzjmRklZsXma3qiEP8UJS4VF6KMJ5FeQsrN0d/lmi5v44c
4US1ZlMrlO6K1aBYQtJyl5TO00R4685G+P+gLSVrKy+OLlVrh2Gd0O4gGlal+qOl
RkAdI/DhE1u2FgqMfMzP5ikDmu192av6NCsbEMNki/TFpiiTo2KsyNKOAvP4jw3D
cugVBTztaoL5xQj4FSVwHjPwPtOUsMMIOlO0ih4oHXlZgrZ6c4HWFHa2QU3UQ6UH
Phsln/NwPcILXSQsjq2N/g6ISjXvQLyjpkXTh72Y28VitOkip61tyuvYvr1lSSQP
TTL99DfRhcDoZ5XXskU3+6NRD0aVIeoxDn1TE2ZZDmQgmPudYqNdw9HauJEwdAiQ
yG9mt6R5XQpva8l1FG0gjEGYaeRcA9+VNaYVigwim5nScJnZyxnKHH4nah1inSi8
9XN2fpjP2MT69015TiC4snpXrtEoVQ63tdb06L+5QSjWQKRgX3XQvG9S5OkTM482
aXEH3vk0v3qy6zSoSJgPfSbRFHqnb8tlzUwZtYCBySKOOigOnx+H2E3j6k8Fv1TX
plsm5B4e/sH5wv94A3RvoXAsj6Ctsd2y4cmgSwut4Nv5eQ9q800A2F8yRJoTPo83
JkTIA7ZJ9Jj1Hf1ziODM21v+b7GpwVmh1iuXEndt3hJzZjI1cgn/QxJbFEijf6p5
06pb6xpgXAUAfkqGzM5eJ+npzC8paAxgs1WmAbNu7H/tVVmuDX4BJjY425YtyzJr
13eNFMGrsPbAgH/rnMbMyrtJe9JWrYhE8un/4hFsBY6su82EN+99mwRQ4oNlQ5CO
NPhZeNQWdLOTMYOsDFciKEi/dEc4+1FhBDNyS3cKTvsAdmKluoVdzEtNZ6li689G
pucNVZuD7z4rCn1ooAe6AOiRSLMO8SzSQSyUflHcGkOd15+Ld2KM2WxpqAmoPgFN
ivsrlJ2eDuzuz1gSC+c1+3bHyT+UqyiE1Dcn0lv/nBxYVYeFFuYqSJPMr7/gK9dO
dHwYLHx7k2KffCLt2PE58JZZtS/Pj6v7rkp9ELSUJCX5EAWD8fHSwNN8zbjNhleG
uliJa5D++TVuT2naQ4ZAoJjHb6MPeMK7ybM+IpllHouYCLubZBBM4ho/qxdQiNy8
ZSTa2h5l2d8bCeH501o7osIL0ESBG2Gq7HKoBfvldXlBRUtyq0ALsF1jYnav6RTj
YM0AD4oDV6X2nu3nonKnDUx20bzPhdCpbfWto+Ge34AlyfYrjX9fL+NtpkWuj0mq
HiJDhihnWeYUCVuGTlYhryfpEDR3UATP0RBXYu0IGXh0/xRhZl8zuC+ocmxxo5sY
MKAmERMZl1qRdqCfuBLR3So8M6bGV2LuLQKicDL2ZAekl9UM6SEOzvuFODOCWck/
xTEnITzSDzA93fTOUS6O4ldf6vbRckj9XrNFbAgGqvQeOqEbzEjYgrlmfCl7Z0RQ
mvbTmLrP7cZfwEhFaZqzGlHYpD209H1/37D5EA8STpC0OTYBSbkEuaRuLs2aSnfP
IdwFO2d7Pmd61ttcGCPyWJbzR0v2fI/NtEF+8mjRj2BJrinXnBKjxjoBtmQ1LYkK
yQ1IOOCrYsEGkp1lV8SiO9fHGiYslRUxaAbxwzdcmAz4XgB6CuFkzeka0Fj5OYQ1
YzG1tyFfSD7ob31QMqTD+caFlbTJj/MY8RGqPUZ4Q8aMXhrpAtgVjIareS1/1haZ
/vWqsheEYenCS8PzuUs9s6w2irkjxUgxzKVMmTQeGKxZ7DdvwefcD/56ogkV0V/Q
aYhti9+GPvRiDdaS01VNDPny1Ip03C3c6q4JbT63QrbJc1heIEG01W3/28jEQKzX
uKnkEDUFPFoxJT8x3sYsijImNe+RjLJ3Wz0fm/wNMo4l41/NrwtviJ1QyC9UFb5d
rys1uh19t7RZXJvMbqJ0xCmacKR8E2u3koC/sTJOI43Jtf2pWwJkcVjn7hrRwvDj
lxZ/upGUQQ65A0zaUGF2RpeXr/9B5HcHwXqCo5Cb+hSwf8eoBuB7lpiyP7i5Mgo/
6AWiMqWPBK9RI7IwkVqdLj19G6XZTXVEkg+tJbnxc2O33IGTjvQB/DnwP8hW5uwB
JF8RR5pe//3gI0LFNSWmGIXLoR1zCokNNegGABSQMj62YwOXYArrrj/tLpj5XieZ
t7nDstW8Fg2eZnZVn+iQH4xuNXlA1vWqU+z4DNilNSZfzQBXHRJIdL2u2ifU16ei
PsAvhaVCmzDq3MkptglkrXhtrGFsYPwnRx3gQoksOuA/jnqO8wBBy1Bplp/8q2Zl
rYeg1BTQAUSTXMv74zZPRdUHhUowJ/piIQ1010lr1N+iHykAsLKHjMkSOsNBVymb
TN8pFkeHTKEzj3Y0xeGmENu0tXln/BdhPkc8P1gKP9d6kAM1l5u8u+5GpUtvIJk0
qxb4d1o6x7IhEoC5iDqkI6T1hCi6Vy/owSA8G2W/YAFgnamW9lwpABK5H7vIfbyD
2bGV8VMcb3FLEsRbR3mDS5O0kmbHDLuRTQVddYmBuZ533dyq0nI4u8pI3x5RLlai
neSjQWwOfKrnodH+GLj8eojkK0eyAX+U86NOdFXwMVg5RFL/P7u5ydtRXyWmDur6
+tkhRQXbnKqefX3gUQm3uZ9EcB5ocrLoSBBc3GIUv1ZX2E2z6Lx0+NqQqnqqkXa6
A3OFg8LZ3bG1EuYYlxqKTC8KyfcATkKPG5/5Ye8Z2rsz8ngM7bNW/CR1e5v9toho
r1lKcwuS60c4LhDN90qm4C9msf8W9PBlDSVU2QE0Db09yKDKGFT3UUvxKC80FxRS
l5oZFcVrYysDh3z0chKzC64W0YOXDzHKyxWUnXm+76r0/AZoHfTXoFi0H/Wl2Loa
BMzO6jplPiSRZzbQFcPnPFhMW/HTz0MzoAaFC1doaNRS1ZWFUp/Qf6SQtYaA5roX
2Jon3+gYV2qE6E0yxhZKL1VmO/YpVNtStScacQZTT4ckcE8AfnyTif4XS1RD2uq2
2/E7jDrPKnS8pMA7DwaUD7fVSWoU45HUudkqQxtvIWBDpgaQrPOmO0DnflfsTgyx
qVymZPv/NrM59KzbNnW6GmQZfb2WEmZ9Nt5xhTK6RgetPKeqJCfg+0nmsenEKBfy
43g+9gdomT2tE473kK++2tFvQonKv5bdcUiWpx14sdlG2stItvxgF+egY+Mn/m9a
uF80ktZ1Hi3izZm/kVHxSnWhDSbSteAChPn3PqGMV5pxrxX/h5DoiSFja3i1g2Uo
oOa2LkxsqYICysSvBTYxsedUbiW8lMHXobRMH/jSlxNM78zhrZ2cggiXCF9mxJK1
z4BblCrfPnfTLuv21kHR5aVV+CHg9/ua/Z58GBhXbGBkDFXLSQIgN2hFvrVt/vec
rgrIC8cOqgFSpq5p1JggiBcNoXIoSdnA7lWyJgCNxjG7H24f2XiFpBClwzGCEmL1
N/hio1vbidlFSzym3s2JOThIjwU0hPwGQa1+AegtphbEohejhbX7tw2qeBvAoNcK
bykWYEMKRP9OUJVBBjpZGq769F50sv++2yflQmYlXjMyCi9fDRk+V+/IWGfebsSz
Z1rmSIjJJI9GrE1WiZGij+bqW1dTy+Y10Dni2h9cSQfqQSaJFcCAdVC6YhMqGObE
oh1R7FdrFJPo8nTuDNyniKD7kmvoUzQX1N2nbTGt0f72bGoaquoq9uNBWg4A81oC
7Tip72qzuSLC++Hh/WFhMi4UaN/i4F8GCjlFKPw7Z0jqHvKouH4QI3cEKnUQyi8a
dhproYGL7I9ooedQTG29i5EK7/nLzltAUlpBkydb4B+cP6Y1qYbbULszrQ5k6UZ5
rVbofS/hlWqwQ2R9wnnncCCdtL4+3a9PyHx7wJToE80VcBl+ir5Eqv4YJvlAxdql
6GBFsreXPCjuxQkuClDmQ4OI1IywPbsqn8mR2K5a2ezDjc7dIH0vpwzixH36+cMp
EWQWP8/LavmBkY4L7rzniYzKx06h3/iyi6CFcod/LkKirsGZMBIAesRwgRbK53Yd
ZqTDCqFpYmZ0sfI3ZDV9s6Bos2yGzg8Tzc8cg35wp3phr/zLzx6Tn6ev7xtmjgTV
e+PZAST3rYzpYYxWKrSKvXDu5H+eyExvKDZI8j5pDfgKUdOvBPuxe35GkMcoX/bw
aSWJJgw3UriN/BX8SzmmYryqn54RQk+IN0VirzE1qlRbZN0YaBLxZprze/qFP5q4
Pfky7fQqXxV5+D1IOnThvpvpiLFOMK2fboXSxKXfR4PNvHrdRapzKxOnMxTNWiqE
2ibZFzdJC3CLeGPiWoKhiuLpJBlHG9fsMpjPYooWsUaS9daalrK4eu802pMZs+on
Tbjo5jKfqvXmA3weLB4LuZ2uCNTMYIEXZFuyeuXKJ7HTq1tPlSDRfZKmmyVd134u
UCa1uiTePiwOP2zOuBZZFns8c6C3L6rIcJUCDP9/kalDROW7SSQkpBC+ZskYi+Bf
PvLNx4T+s+Cee4ruFRQSYOKoYnrGtszMLsmMbVvwBLueCWczSsh6nc2bG5NviiKH
IcaYCh33BnXsUJfP+MsA5vUbilno427ERVTPbC5+c511LD3VNwpqfmwZfjyKnGa0
/6NvKYQ3S1E0+UHu9S8inpkYTDI9qHbLnUQEwYJZZEtS/HcbQUxuj5nNGWnNjfxW
6UXpClZvgfd5KvdDFAzMCBlxNmYqF3MO/R7lgi8fhs6mjSNO6CHvkcGEHC3Da+dm
eODhFgh9CiacWlCdouL6NeAS2+oU3lGDRTjMx2rVeOH6FyHnydHpssUEtmbdm+Rz
G4JvURhKWzO+hJD4EZvJj17d536FnhMSNRyZOnWbeACHcySqeG7jDQ+2TqAbLLM8
BMvYNVxCIxirpgRz7SJqtj/PFvNrL68OckTHXH7DczCCkJHqoUXUmaivwPiEd1d6
DetnoV59sQAKR7HZQbw2UEwqlRJto3I+r7YWUZvnf2R46hoDDGa0GNekqs4JP4u/
xjCK3lbj9VVT0gE9ZPOVBqBaMw3j/VPu6RGM8e/S9VsC3r6jpvaxlkEGWbEpXUAM
h5Y/XmfPHSUuyb7G6dj0f+Ed5nQ7C6FQTdpwTEiEskaPJSkV7QRA+xGeRwToCECO
hYdYvA2Xig5g0/H21/knfC6MGTDyM7t1YVvc0BEU3GxFuMhh5Sidl7sezNYsubf3
t0Q+px/9+HYN+uZLcCf0GOplnfTRLpCa+LMVbfqImyf4dFZ69U7xcIzAcUPEWIKL
Z/gwecMGi4523xfflFMtYSoqKRx//giC4tSmyr1ll7PHJtIQHA4qGX9DxBCATU6g
DqDoox6NhNUIXkFyGFajmcwoQ6Mnoi+JCk6ncl/Rwbicp8aaMT6+qeQtIjFJV/Hx
9XaSOFmCSxXTtqGMvl2AmRfxz4+chH4g1hF3uFksUhiRHuKNCfw7dO4JG0AvrniQ
Aq9dkWRgXGLYGZpTOR3sd4OMUbJX/vog+RDGE0g4Nrk9r0lpD0qh0YbFbgzru1hw
VgBB2wxUi2c5ijH234hd1L4o0HMb0QH/PkugJ28GmiZebfs8sJ79ERRtmVnConBY
lL4Za1x4CJ6hewJwOd+7MnxP7hLaeLfWCLQD/bTlrAtolWh936sMhAmack5v/Bn2
2QegZ9xl4qlVTUt/pWwmONNtb7OuzYboQU6xHUAlwOfdlrTwhjHPTA4dp01X5kcb
ozO0euuCA3sVD8qviZwvBqUUt7rE0Rp+gd6dgXSjRxjcuerfkvsFxw4F+4QLKvSr
agTBxfshYPjiU+w4jAv4rNrMyXdYPvSKE7WuXW2+m9og+DrVKZIONEy51o/yX447
IEB3YXOG8uCiZCjuw3x/MUsmW++KLZDxMbRVy21NPjeUwPFwtMM/6NWIjOOObRx9
KshIlXTBkRuJ426E/uUogB3Zwp8LQKSbmt0EWYwOoDZqcyVLfCN+0uroN7cbSREV
5tfkzHXp9HrFSpQB80rHdzehrDUh1Z8QFoaBSQJArRrGNToRqPNucY4fWNmmUhCI
HWD9sC5Xd4PCx+BwufD7ebjuGfrchOZWEIsW8HgeS8nvb6q894KRmx3lYiobvZT9
ightCjsey6TzQLYFr2CewXDYqX879cj+O7uTi9pSUA0/YXGPjyuzc8okruPS/5cz
QHNQm37PMAS91yHxfy88Cx78qS/r6YO5//eId7M0MS3ejqtA2epDPX+TEBhslrb7
xxJwNw9cOvbY5vcGw5zG6QYgHdwSZYLjQOIsCiJgO4NDrXIzDr80fDynK9vo87qa
D9pjVmwd/u3mnIaO7jargZJIHBJJnO8p1n7t56UrGJDYwREBhmtoz1qVfA56I13R
q7nkiBKeaUWqHXrqbSWifWinkTTuvFxaKGsrinWJxnHNFkPLyJll4De2cdRHVtZk
np1bq1WiJP3lCpuM3+dl+izhiIAM+dLF93YjxIqzCemBQR0OU4hdisAq0hQdK2Zf
VyN7eiOn/EyGEa54aFC5yoG6m6yh6Y0BLMGS/cuT7YZbbhYRAa0d76Zf/OuJ9dEM
2fquGRk9nyvRJLNnXq4JS49k/Tt3bC11+WkVNLb5NcApnGZLWccNPav83JmaMm+B
elYWFxkEgkGCNAgK4d/hoIOC9z79TGKMOfYiVr158w14Brn/atcMYyvoDUKqheMs
K+KMJciiDTByp5+38Gfz75jUht8UeDy99RfWC/sI8uAJ71dmgl7rgwkr7hN/8cEn
pm2HdvqVhd+A9jupAVqJp3L2hhU6sCageLZ1FfkBgW+ArsPoiXOAu+Liy3lA2+aD
5/Ym8GQ8Z0svzLuxZWwnt+pt6lPBJ+1l3d6ZIIJBwaMXECzlKZBdOn1dxdmhDBFZ
HdCiw3XlhAVXWWOQL1sPrTKnL39zhcaR52sC9EMxJlA9N3i7aFu5dQcmO9srASDM
/qb7N0lQFvM+OKKf+LB7QehomELCguUsloxaG1eKqWhT9ljsTkNXz8b9suJ3NQnD
Zv0sfu/kICxingmNvfo5PLCaNvOYZPp/H0rDOVYO8mWv3L75Li59mnzQ7VLGpkyO
7ItCnDlyB9T+b0PWDj1+tJUiYoyUGzrmbsi4TqIhnqoUEzkli5dZ9dmUI0NGGC4+
3/6KsziMzSFeQC6Xe46WQTmqB2JNRaEUM3LcWQjp5LauYYH6yezoXMO26jD8+HCZ
u0KpiPB92kfdWLQAC6hx/pruLo+MDx5YzaGoN1GcAMWCLrgmI2pN+G8WNaPc5mpK
T8gUELXlCgZi2pwktmlNQFEbIKIzz1rJvcRZqMu3igR0iSTLXxYp+giKJ2+8psRE
39JGyCmaJp4NWxHjgDKRc7r0InFiJrNqj6pGtqk3foFrNgVxSD+AOwujQwKXW5mm
ZYocy9CyYTHrNbR0X7FRtfdfXJ4wewgEmo/Ol7QZLUIMXYPLeSKfq7IoQds6Ox6Y
bmMuAC+3dMd5D3efeB5P15A4orR/kahqZf6laQJAiHXzmSsc8OvQfYmOq1QReySP
fytisQju751fD04ZQp2bwjaSCOceNVdcA7rNT1qPvzfozU+Rc2rkIsR3TfVSd5ew
IGtojcUYFbHiNkwTwNwhlTLMsOd8jzs/4qdRG2FuhMWEECU5Inkavb+Bl8Oc4YdU
Gcek1AgiYmRZFJxFgxcGXWgYHG3UbcYgYkqjWDKebxZXs7sd0MHHPIC3DwTwR8Q4
exWemJcIc5gqseAFkXNAu6FHyyKPdoaZCgGbyqHTGBc4mtc1aB77L6kkK6i5Zc7W
NnaiYZJ+Ub/wWUCggR8nbXMQlt6RhBn388BllvDmD1irxtfdgGvyA4kzHnG1vkIb
VOmdtNdn3KO54TSnErUbAXXo29bN9lVjPCV9AIKw/uIaYa+MZD/OxIaV+t6sEDZ2
tTJ5T9h6X3s3Y30vjKZIkA3IcJH9DqMoOh36e+3gOt0dmbtsRLUd8DUM3APZ82/f
X4Jwt3119M2AKei69VZnpsqOAznPercRolRE74Ovcyhu2yHVp/LdoHTkG+vqBqqN
pP5FpFTTCIegaV/Eex+A7qBTh7dcmgNDaKeT7AZoYoXXjvImtJMiWUtKDS8+DVsg
uZpkg4v6OWco1ziEe1DK2plzxoGjBowqxjAG+LIkPjJPVT3osV1zFQk0EX9EyhsO
Hd0WzDnnh6qzE70zLiC4753CQ3YFhWWZIen+ZsJWPvEsh0smZ1mEmDPYDp2mlxXB
63xgppHeHRS8gW9lV81cLUUHU5UWkgN63YRuLzExpkgX02OZql6FPI8+DJQnmg9z
4KNAPMC/9xW7XhoOUtnU8og2MrqEELkKAiPc+fZn8/Zq9yB8/Ep3h4ABHUwpdI4B
o8rs9i5ch++rOYy4J6cPlmzCAvaSHc66V+gwHapszP0r/1igHQped9TtTLND+Pir
9noFVjCNWipbdn1vgNf98lBgd9Ftc8qBv5m1VmFXeAH8rv9vWNNETyTd6fHLKgYD
zXNqOT6+fc38c0nSbBKAMbecHr3OZkwU6mtVqm8wxuAf6fAF+mVZOC8CqnpXYg1y
W4Y4PK/tr6+e5Ed+QiupnnbOUR48LtR/dXEYMyrhrfFKTHwS2NH01tn/XMR6xNkh
OuxQD5gF0H/ZvhSWZl13LHz08KNqEKGvQq+KP6DKT4Pllanbdo8UDJET1mMCP5X2
Rrey+VofQL66N3CvOQxTfzp7PeZQ5YeGWvxQCX0EcYj1kPSfeqGV7aR1mCPYwOHn
ejeFBXnmHMoPjtBmQGCmH01hJnR7B0HY18czJmMzYz1qqr7G6uNIg+to2N4dFkkA
CwoCEM9EABbo46B1tnGTS3cSmZv9fpaHH8Mu3al2hkeRbgVeZso4Xm7+OqCDX9lv
5Az5dkxjIdC5sk2dcIQriFYAqXe2+ITFHt8zAeNxZMUiykcVICaheFWPdxPXBzH+
oiGcJjPUGFzT2G24MZc7TA+oWcsia4yM+j+dhB/qL0pg0PkWPZqYfy4dXk9Zu4GS
ylOn9+ve9s8o60rb46oGuk8EoI2AzSGz4XTOQzZiEvbhx5wVrnkvYSHzV5nu9nxf
3o/e+59dO7/ls6c4nRk8Cw1ofG6UDcLZxJ9HZntB30ho5H8KNLO8mRWpN4AvNdD4
Gyb+9rpLJOhZbbmX2dMGN+lGob5hOHisjfOqqeYAvPjguOoAbpSZckaWIrL9xVyM
z+cgX32MyUm8ZxFe6aba2fdO63Qg03iiwEBjNV4q+yvsrzicqXpPDXX/pbiZROwJ
J3Htu/2bmwLUf7pPHG88LJkiaKZN3cNqAyP3Gz6607YYo69Kukt9MWMBHR10Wv1M
vMycckHXo1/SI7o7MYo23lutqUfHBC5Ui5KYT5MysI4wdr2toiz7NzW37RyIkrrB
g2B/iy5Q91xwUK+LF1acOTnqYdH+PJKNmDQiDmNuOB79ybBpH53Q1CiiyrI4IjqY
IieNUoTvSzLMSHv9fiMM/flOKx2XXKhH3sPCBJSXy9nm0R1GHGVA2eOGxyDfUIji
BN8qx5AOQthCUcXgQc6YyisHISykWQ9u9VDz/qG2pSC4MvG0i1Ocf6mUFw3zg//q
7ZHycCmdV3MGe7wU1tJ2wPA70hdca8TVl/Ru0dZN95vxKWvcTgpWxK0kmrhTq6QL
D5tFzZbYwfvfecZzX5W4Cwf7TnLhDFyUoJ1UcXnaLht+8U3ERYFm8unSPNMgn7/D
B3sJM1XIOS0n2juxl4oD6dqCDRrWQqeHwFusyUrVf8QeLxfpvtfWq4nYmTzyH9cG
Bjyk7400cgT1xirpyEZDsZek94tR39ObEU4izIyEMSXx4NUwbzCrOTIwdsDeMRVb
5jn3z0mRLDyljppcd0ONgVmQogsyMF6HUxFKGwr3pNBfgzQ0a8LjpojEawc1XNBk
vUnZnyDCqP9djaiKtWXz4rHDCXGHNrR4gn/L3loEw6xQRsRAK/IiHOe9LG/GHmgf
CEGtTRCULfgpeJwGbNjME1aiPMuVG3cXiCpJuorMW93ZiuU91Lc8NjJx4bNOmCX5
QE2fqitMl33RnMibvowiP8qXuq1yXVNl3fxp7FQpi5e977azsJSSLdhFYLzAK6Sk
KbArsv1UObd6i8XlwEmemmQBLjcM3R9Fttnd2DigGlcZfi3hE4yKV1/8pvL1bDin
W9R85l+WEbieDVZCYIKlsXonmqfZJ+gqv3rtSahhrqHMeKYM+Dmm8DJypCH1LgmV
CdbYUMdVJLjCkb6A9H+2Q8AR91MXVFeoHNGbBWKbQ7DiCVQdgsWKUrQaiazW20jZ
HJKrMywCN25da7IT4YvJFYRvmQ0urbzUeM+Acy4aXN79WPlOhvNdHJ80I7MHK05p
t6sdvn8eyUIvYeyMDS2auMdNCGp4PAe+yl2LAtPAObKcFI2HJxX+bwBTwQRY3iv9
MHOV7hvSN2jPLm338onfIGwfN2JTrOlY6jPdCk7QA1UGm7AoI5Eg/BSF/T7+u0Uy
BoQr70zeEJlB4JXY+LPVzkzZ9IZX0N9O7kY8yLIPRYsQNomueU4HaUowxdyNFXO6
EUsljF6hKbtht7LbHvznZxfTg/Xc0jVW7T7EBFN0nRywyGDyugRXhZ2uIQmqdviU
4ZTQEBN+xtGEA+a6txBNkDQdXAffd8qwCcoBswoeg7AGrS6ktdNFI+X7TWZv9vIx
D7KxMnlXlGqX1py7sJguvuBLQZ+RGkBYbtPeZ0hzPUIyDXzm72TIL4afCblvWCoB
DZ0Tg2SFiBlLmTMmqQCFupUnRsofEPUAgW4cP8hDR85LUVIPWpyEnTRwjhTkpZQh
AZqDEvmCsATU6VntCfBf8AWADZYFZVGb0uNTqrKq2Kug+UU1w+5v+W74icOmCnJq
91zXJW3oZlCfnSc/ZCGz0/rMYY0iF51DxdTee+MJk2ODuyLrVRPURQDrQOcovt+S
5ibT2jVaC7tAnu6Z+rw7nz5Pzd9O90s5pEfbSCvLwbL+uHyFr+lUXqFMRoKgdj+z
yeG6uA260+JtauQt8WkTaIYokDtcmRUcLz8o9mmeApsSEliuM82GLnhImcFEfaww
/fzo8/zAMANignYWvOM8ytn94cDSuOGm8X9HuaVtEmnfXRS8/bg195r5UwymlMs7
TLNApD2TN2ZmLaVI96MOZXp4lpdO60MnZx08yCrUv5jntAHHvNMuU9jfWYbTFDDe
MzaeLRz+Fvp+TcfVHirQDs54zRlKYhntW/p+SBVk1CpjJZnI+JDQMaFGJUGRWTG5
YjWHLbTDd9aB9x0HCGSS4KoU8L+Gyy2QPH6nkzRjG5+9jkLUyft/XTcP2TF/5fVP
xCmTjT3c4LS+wZixUKDv8FgdsMUmWPlTPeOTUKe7JX7zzh+cZE+aZsg4ivShHwpN
VGEDXFKgt+9ai9wyKJhdP0MfE2MBqP2oQaPvFhy12oEStBrB9fqwOspmezE+KxIR
KhcqCrn0loRgcd2VMSGCWfszS0WD2rPuv3BsTUU1omE6T352eSqrPLesHYqXLrKA
BI2DPtrouJ1CeE4X/LLdxRUYhdyDPYQqA/KGEq9lLdAchQ/GSkbOkxXRFG6TQWPN
G4TWET0uVCEvTdqh/Pnc+Zgw0MxUhG/l/djtb20GQg73oYknbTNCfc6YlTBpyreN
VbzdqzoXsopBQqrRrbhsheB3KpCuYP+uzi15AuN/rVR58zhnw6uWdibMRjQQRdRn
Rhle4UvXyP7CrfXM0M9WGSxdnVGjzASDDoqmGfQMloOqAZV9N26DCtfxgg0xRnpF
9Lyx3rX8t9Ia9nN77g8xt7EO33gSbAJqMwAAInSzvxjGa37lIsgWNyAu411MbsGE
SlaEDzjuXwYThY19jC/L/wZz03wViukgXwPxy1aXabJLBAi/YqaRbLCHg86Vg6oX
4qiamJ1UVoOBiiGj4gYD2oknBo2LGnFz8h8bWtnN7ECedqFxaHfxMdopi/SbNr6a
vkTcYTJ3vfxyMQDFPW3LmJs24+nEbUrDUktY8rfevC1nnfEHNrM/8ogWT7Aue+MD
Ll8S+rL1Vs/9lAF7rqktT99QTBJAeisvix0a+AOBQLwMu+y+3qFbSERf4TD6Iowt
+9bJXK6LVHKsgvxPRsn014dkX0SVr726ine5aEz6u1zBdRQZiGK+YTQTlvbN9geJ
zcpS5+kQwKoSqRIH11zWI4t+6WPC8zbAp2bLGY2wrQIPS4sNA3Dt/JJfN4TSIT+t
1vyoDB9pmTNEaPHaBetXLjzEG/QMEoi1NMP7qiG+Bhr57eEoDqmRIBdLTnMM48ph
Ppcbg2BnTVycsgmVpMc0a99Nf1YissisATc7hQpz48HlUCm6ghcYkCEwyR9xQUtu
ykNAcpPN2CfqivB3mB43rDBQmlk79nlLI1p+DfSgfPdT3l63N8U0LIKQbu8PdFaj
A9zxp97MdqPy0baY0gFbe2k1lIW2OHkpU8dOvjQK6VgCaubu289moa3w/sKPfvgk
M+pje7mkjXY10pJIYSO719PFVd/y2HIMpm9XwsKo8Hvlqv1i0Ifio7/NznjNeNTz
LeipxzPf1DSwgYDf3+qOWg2yjFP5PsMc5BTr9ML3IYdHhg7epbtel51ZRyWcI+pU
cCSxJKzsO7mA07wWEGk6vghL93sKvJ+d/z12dEgHizlFuc5nQ9OT2SEoEj0d/Q4R
42tgawnLRXfQIeNb2I8/f+uzHvSepC4g2lX7z+2qLojeMUo4CbIcIyvMRoUuNAm1
0eoD3Owoatg6q9+ALr7vzzX78D9ywKYQJl9GY5Gq/WnFQBgqbVbStFZewm4sk0jL
la88qgACKUdjT8ma8AhUn9Cjv0MUPhqLtW9Eox0wO8PD9/nXfZdmCl9GfB+OPnHd
PtcE1NMnxUQ0+NsaiaGgWhlei1rWJ2Fvrp6zwyD+TvfGdFE4WjVjbdkYJHyQSI5Z
hJDSr7ZfZT4Qa9S1hKupKVenUZ8Hq6BYrmOeEiRW70Z064sHhgZvJBfqQSnbhhcc
AhjnmX9koz1zenZW/c8+yH0nUkAuIsGxQK8RaVtaTTpazsz+Ml3wZX5wPK2+4/1X
nP97PQefoIcVjxe1hRuIthmVDxDfK1HweUF59jTEH2iQT3TDlP7+GUo5I94GgiJM
7i5lVjXEfIrK5JxGfsfzK4MboffR1HX/6xbMIGcQGT/5iR2t2iC0n0O/mM6P+2lw
oF3a6qsI5I1YmqHfzIVQeHiRWUaD/Xm+1NYzaDEbgPaMReuFBEcAkN/yR5PibWnO
VVohR+hWUrJHoNXu0LpJaVZmkxNiP0hLyOnIs5hxttT+ErhHB8GOA+6/OnG+NnuH
HboYSl5m755/A+m3/T9PkPNzdz+oee9oJVo+2eIeWlTGQgKQg2vbLKGZLNMJgOwh
yudrVAhtwbmKfzodnBHpdAb+Chjw7tXmUAh3RMDJizRiBzYGlMvD/7C/Y/x8fvBM
EjJz4X5sp7gfcprn3oLeucv+xiUazE3WwE+j8Zs9bay7xL9fItRE1Qgs0JknBGB5
KEkSX9zxsVdT/mFcXo4f3I+gSLn9v7NZHCYyRd4nUpfpdLNf2RwsSDNsb/OXq1Ys
GuogS3Ok+anVArj+f9og7giujuj7DaN/I2TR5hPluZ1boJXKo7EEwbVC9Xfk/CKT
hVbzg8XmCroxK+4abAR3F4XDokCOmBNRxAi7zqTxufZZSWYWod1htSF2e2k6jlIb
mkiQr+qnNQa4grTFQ/3/7bEI5GSbIjIIP7ogP2Efw3EGw2464lA+mCmQQLqr/RJ9
9zYs2ovZNkXhDyxs3ALlPVqwe/MvdFgtsCiKvOFaiq87c0JnmUD+kUf7l+38FpyW
KtaFEBdasrWpGAb121XNUQzb3u3Jusf1ACODhIwVkzo4rzd+xiRs3QjhI6cA7BzB
cNYHjJXjNdlNCBrvjgQqnQkSoFNyR5zh776iZRIvOWXt/ujvqP6BiHqqb2nzuSlj
h9DskPhP/VTIOvAIquQcrAenxUnv7UEKb9w7oqDW8u8YHpjr/utx7qlc2/cR7Ige
3saw+oLV+Zox/jdoXKHLjMQD0In96j97sR78U+NF02q0w3nOzyEnQxdyf8KX/78U
oY+CZ2oAOtKQZNdcMuE6/m42NDvYpDrVjy01X/NwpMvt04vUIyWetGBer4oVMbqQ
qAG5tmGChIISY9/8MoF/4DXTMtdEvmEG3kTNWseW8Wm8VfBe54LEZ+EKpmsvioxl
BRpGItKN25+LJn1eeygts2CnzGfrRKewXFWB9SBAzn4/vMfZoXIg5rFBAcrX9KfZ
+1ZqZ52phP5ByRtlyFRssdQbrqfh+oxAMH9JAFdUMeEXXzJlr7Gf7vS358vNw+z/
9y35eBYcplY9GyEuQttLDxtw+WZQ7WMGIeBcjUlRq7ImM7v7FS01yQQK7SXxW6fi
IRb3pVWeYyDNssSL67366y5uEaeIdbQ+TxR3VMpUfs6oUd0YhhSZONtABwwbp8Xq
QHTTsZM1JqVKzGBzORBsgsChy+MjSseSvpEa/A+ut9Lw7b1IO3yEhQEwlyiotG+k
hZZPuac6NlFKmMTucclXqLPwETWo4cu2eYu7ZtkTe2zr4l5EI24dXk9g/VumthXG
3E7I3wOKqeVsuXfgUCsccKRmZjDXIRoICPAv3Vj1AKnUzZ+EyXpKqxtxqJR/w783
3x1sfGwckxaPNew8t/KJVY3WDuua44hrAJzmsJxAuVPs2GLW+JZjkwcUe1BJe/pn
6/mDzwSsvcp2afJv4JRzOTjYGbV+DRcuwNk8CoNcXbPQbbIj3N/llUu8U58vcJhn
0yBk087mAIODQ2eF2FeeNXdSYa102QkYTqCTlAMxlbtJhBVT5eeCUGJh1z2/49Qr
JlVe25JbfvKNmVB0tVfmASSsN7U3gIL+LB7p+YW+BZ9SblTOssXWhMZRiV90lGGH
ot4/U69Q+7vfdLuYnafM9/SkgeO6ZHv/ChaHvUHgnY4KnExRCej1fCAjKNFIN13U
/EjMBCBvTFIRSRWFmBe24s5725No2HA5C4cRX1+bJJyXHbuor8ElgyJHckpnXwwj
y1h7KyS5zoHGUWyq2BrGRVX8+oi5HiGVO9AeQTWtq62enaSQDuCUPGnGbeXqU0Ah
4sHonLo1oUUm5PweJDVeCdCcLbKXhQ4i428er3QDhget7oJG3ik+MZBYoSP2BeGy
1l1u4i0nisgMoU6R5eH5DBhUKRmo4x2GlFICWbaWTmxSZAEFqOhmbEXccV9pDDtb
nUajpj1UKQcF4j/GSFluWH8o1rdU27ddQ8iqsuwntfLP5LA22S04WrEXiLfXn/5X
VGrpMBvdNCm3g+W1IQEap19pt2X3B3UyD46q1Qo7DKXS64omamKQ0CM8IZwJueyf
cfd4gatckcF7OT8/JdzjreHzGBv8eVkk8xtWAuRgjVC/P5YXt9+orp0Y8RDzbSqb
CCqZboaOcgjoNLq3h7Eks033IwZuW2fqAtllT/Aa/pVi8nOuEnDsYck3GHTp6SDC
HYZdlYV7BFgFyC07HHSh4nlfbVFjv/wP68yid/kDivnOgi2oKmlZ44n2Um8Aj3PJ
HHyv6egMXsTP2zvZj4SHW2MKh8syqufdlaYW9g3sWzv0x+31EYnyj2kVw+/X3jGz
4TM9mXraOD9oogryL8UcNEcFhVQEHksa68OMLFbjHfH8j/Wuj1Wsu96Mf+4h5pjx
dDwR9qrUYvdb/ulENq3TBJ28XTmrYFqpXuX2/olqV/TrygofrMxvxT2KMp7WgAC1
Rn3XZjJEFcR6awMmr2/OXwA6u2AsgAYWyRyFsEKifp5cCEyoaLlgNbjMYXsv8HFh
g61xtEjYIiU+N4O7Xy6sjcUVS9puHc6DEvDdwQH/zRnHDhOSuVpV4wbtyXmZpPO5
xlXqTO7qW0KqYHfK+TYjxhQM67hutkf0p8yYyLoq4ts4zoP6PZDQ3ZHFouB5tvnF
qN71ZNuXF8DVpbmpVCJYUm+V0LeN4hj7B50mOj5M3mtxPG4D46GToQFWIX3kjFiJ
6acxGg0lFZy8xrxjK+ekN7ItHFe7WrHszZF9+sX/9Uy7blCuFAYh1K8HvDixqSU5
7G9wLnIWuqatk2qcE1ZVqfCpxpM0BtaZ7ljsjELouyKUOgdW8PntIvO12gGHdk0P
2gCyXExwzqEIutauLKenpVMRgUm87278WT920tK9rUy8e6M5YqL/pZ+0W8lz0ipO
KNDTkofAgJ798XGDpchB++OYroMwVqpCzUmYcmv4rubLUGC+wrwPCJ4LmWKdPyol
E4IzPjhqERhWANzLRF8YQSvrbk3lnj81CSNDjstBcFXAZ+Obnu5m+x9nI0c0uVcf
ILgGA2+ljca7r63/4Gq/7BSQFcZJ+iJUMnwo6DvfFINxulZ9qguMKmwVAO6ogBCO
EfYY37w7OJjTSfjua2pu4ZMTMgQDyAc+W/QDSVO+subrBnP0nCI43vwNqynBFGPC
B7IcmAg1rKRjmbUFMyYJPeaNv8oFawV50pSGyD59HDCIHaDK2uSr1y9C8sT8d1SV
LQV7AnPImqz4XKMSuTIogNWfIKACfMEEL45Qb84zxejcABaoTlAXWfrYTcet3CMD
8VEbF/KhMuZBnbNpTVCSZ/n+aCXsZB9F8KHl+YpvcR8oA4j+E/hV+DIxljixeGQX
c1JjtWmbDIYbkEf33p6fYxF7D0PbHJ6m0WICJr4tGde8GscbY3c9yNu5E1D5IV8G
kdD++f47zFsoH+8EnjvIDW9SFqE4oqgnj9vZj/DhVITpznZDgOTqf9A+5IZIYPSd
iPdFUOcA7FvHOP62hfFSNSyIsdsu+2fltGG5St7+WCcE3a+s50ebrXwSz4Gq6TXS
Z/Gp5TFXPwqN9RodqkCW0Dv/UMDguAqaGyAzA7xLhKY0ezMuSLml7P9cQkIJs/VF
uMBgK9OKPi8oY/ZKumKuP39ulbnJ244SSEkcveKidhn4LftUKXJOBnwUVZwPyeCD
xPjHfbz4cx624D+AgxjTqCDiA6CHBUh6yrqCFEg88V3RKh4fgoW1E6cJJOdrePAv
M4yKvH7va39ND4QxrOZoQL8FtuCWRO+EZmEiOENF79lpPl3nrVh9rYSDGJhBSuVi
lEQ3CMuMn1O8/nCg1GB/xUqqB+bFFImmHanvMBSZAdVuNSHA/htUmOwHhor3/oh3
5ZswlJvAak9EqYXQA4HNjayzJl/tvcHsu1yLBSnIVGG/uobKymLuux5nke3413Qp
CV0C5Sfn5PdKx3yFHrP84l8M9G8qEFJhvOb1s2ddNbiUvDapcxxfHhYJ+ZLG34Ml
ZmRtfh/qwDSqv2vl31U1EMa93pbsIGILqpdgQFGCRkn1CsRF0XQVb0We8aASMPq8
AcEI5mSzDbxcbZvDpUlQNIqPpjPXKW0nvp0hy46nSRXP8Sl1BsNVZxpIU3Es9SDX
AdUV5JFtzH0wUlrPFS6reMob8Ir89ITNzcSX5hBOrY9sHv3WTMdcpM9lXghvRv/S
gXi10h+JG9XC/euiJhnwguhHPDL+pwgSWXXaaUmgoyTEQyNKqtUAZRlTjLRx0NZc
r4RzGFo/dQl6JKBLo6w5PwA7RAXufOji9+APvLLtRjdUT+5K4i5YET2ejcIcb9BU
+kntTp4VyYcsyxADZdhxZ1M1BqKx2mWIOZrtU/p8uZAz+SdN64ahpzUWVeO56yBU
tioM/qNKyqqWebfv0v7SJLnKGCFanQyshBBulEnA/XLCEv5GbDyrFIqoNTSF3UZV
FQd8L7yUFyfqTqEfQ2AYjlEdvlX8E4fS8Nlgg0R0c+kecm0to147IJV80nbq1owi
IO0rKUlCag6mI+Z7bCBMVrrfiUsCVCSu4OihTnkMvIDhLx/hlqjxQd/ftr8DGYF2
1mMA12ckl7lz1nYdPX/raRRhxIskn7bdNsoQRrSyoONt5gkNK2YfeI5MKwqypInu
pyKGeYJa4jsnMvsn4ATbvISCruGZZmFHiZnGmdYp4phQOf0/oTxx5bkdd2CIpAGD
DkJwkCt6u6+3yqtq3tUsmdiP63sfArb7vrwxG3z+/8QJw0GdBbsrXnSdmKyyaJAI
MLnWF4j0IiVXHkrubl9JpUvNmElvTD1SuW0+vFe9sWDyaHi0ZczBwbY99FyXbu4D
iCSFg9SYbiLKSJyPdlAPz1wHvVzmwF6AMCmrbtcokF9LscxrXQQ0CLWzrlcDn0i7
6aU+G5cEzDSfO8mGKTWsqExccd3XAOtA5g+OZkBuO7ubReibhpQlzjVbmuUk2RuN
0Av4/+T+Jut2w51PNgwlL1XPTCyyzOm2sxUOq7gnltjOJcTMTnaquBGLjdxivZd5
VknhqnSj/XF7H9XcQmhpDj5gKmPw8y/zZLUIl76PGpW9YVZBqe9I0RSqY3HpwZqw
jiHy9W+gzcUFTsFozCsBzWmTjAKyBXduTGAhaZYki1jzo3ei0mubITQf+ZEmvRrC
6DiBrlMldvji2Z6mNlQE4pJmGvJ4PwM+AmVkEq7T7Ww5+4dnlf3G8tvXsc3KLSW/
vxYzMyWXb6NdJIHFQIn2DQ60uMhStUUQGPHdlm8sEXxSbuvFSelpm8mayuqceVcn
xTuzbwWCaOaUF7wgKXg1XSvBGql9fOf8KMWx8uJsI9wyZLHIAb8ydTQJdV5F7k8H
2hMNUCoilxTdq7u5SKA1LsQwqU1a00tmDA3FS9TG7+f85B5L3i95MJ7pvi6r3SuD
rqN0QUv+RrXlLkNsWKTLSVk5qJOlJ0Tsh/jl/tyh5j9onnfU4ZcdUCaj/p62r7A4
9RQb1m835zJIVwTCTa0namCHqLgDmWQ7cIh4cmZSrDon1pB3iukwvpO3yrhbJNhv
DphHwzxZs55qT52/l2cWIJDgygqiakY3K2aLaApAxGMqeJIkSdmF/IONS9mnhNhP
jNNXnDN1/+skE8fBb1EW68FNxyweoYMTCFfJx016VVZQiq7Ht9tFevmDnOagfVLT
T7yLuO22XQbG7uOYCG/JFGsA4PPd2tLy2FPfj5gbu6L+Ukl4+8R+3bJWQEX+5xDr
o0z2ZeCtPXbxyVeMLsK7IGQ/2n6yJSRekmH10z0cekt5UtsgDAWAoSDPowiT3p8i
cBT9NRrmctzZLZ5OERFisDalEgoGtmtyOMHOdPWhDR7Xwbio5n6J4jFFMfj4tM5Z
a0ujXbL/946KFK4rneErvXLU7yeaDPo14j0NTSyQbv7ixs9ovwdQhDc2shHIrgXL
HPaIEf99XSlmCvxxTim/OxoCEUz1sxNllIQxfNuA1FzVLpXBAZXAZa+rz+BxUuuv
YCpO+AiTr3nBW2gLSAKYxONC1vO6ZnOLZCuImhf+JSrwTrsv2aWw3CpWSEBHiwWj
lgFfMOhP1RLumzvm94DNwRtI9uqrbNiMD33CcIQCQrvcWiZWyRV+tp5UQ3F8ItTi
Mi9QCYNMMTsG2LsjLWkK811/5Ykbs9PxubHiun4b9XomMg6RHmQzUv1iVT6vPaIf
Rm7+97S/OjyQlCJTqi1/y6tI8SYyyb0XZOEHvQPepF2lqw685gelF/hN8SiCvyx6
qazotUe+EyvJv7xyHcTDNoVhyYbnsDhtx4LAzShfuIm5uZ8w4x6t214jtog85nWL
iW0Y1XLqWKrcRG96cS0dH7zpiDqqHzE498/hcICpyn+ZzOKZ3KZXPPtojNAXU1LA
10Nt2jBo7okdNhSRlynx3FZF3Quk59EA8rg86vN7ItyZ7fdh4U3Z2D6Cq5rNviW6
mPcEqGnmejldAmewxaAti1gghMvh6mkr6jcHf8Y9sDYcZTm5mXLnQkMF4ppOUKVK
4hatu1uqzHQW51p/Jp+hRcTNU++3G4r1h67znCj3rccC2Rm24BhvFMKLXcFTatRn
AZmrS8lovtuCzpxJovkBLEFnsdUpsF3rewZMTx53sMKSLtJQziY95YMkdV/evDi+
pain0uDAmpbzC7Kw4TvMs2TktHHNzE8nfxQ98JqaN86eYGiStSOrxmcFFnVPBDIR
UBYWyUfX4YulehOycH5gHGQ5G4ftYJrGUzloCmwgAP9V6XLFWyDfHZRvQQM2pMFm
j93Vmmaxp9jkigGBZY0VP+PnJ9MnjdACTlFHEhJMuNHj8MFfOPoiW5bFLfdBO6+J
y6pCSGAFajYcWfJlTJ94OBxG5/jxYTrntEAZm2RriS70VtxyYpr3xgUDzSdNcuXY
RT4HuqFVszYdoNeF1kB1xKuWTXCXeio3+Up1ZzZFOlNhndN/cYiCuv8Y1SxOKkih
5e3rBT9mT/mDQepvAnCZ3xe/oVAfIE9OEAFk0/fpghodTCv5Iziws3Iw601/LuMK
pPLf8PuO1SJ9xsc8uSZoj+XTdDQmftfKwr2/PLkGuaP5zxZl7v3I2jeEv4re+qAi
AN+7KhjKPxBexbRD4bbkoxD7nwzxXb1pZyHyJIMg++DYX7h6am9L01thw7KkeKgr
6sTNyWPIx84CyyuAksBBQQ1BjQzUnTre6DoA4Eb3NSr/G63X5A3drhtbbq6F6/ez
T/uPG7BgF48S50RG4XGylvrOwqJ6kvbH8rsU1RBr1vksDHX0nKW6wZf4tEEPOUwD
S7R/r1O+Y95z/gfZMNCu8FYzz4rDDR5hLI3WqEaGw6fJfYZIMg5P9asgQ820yUMK
wutI8AO1YJ0fXe3IZtJL9/FF8HW149K4RS189O9vAzCaL7mYWRqv//xTpAN9r0K8
3+rKLg8BX9iahaU5Wt77f2I7ymtw/CL2Zk+2ud7iNVPcZGGeYLepTctSX/ihJgnd
urDa48RmPjManatsjYEbJ0lB9SnjPdxmh1v7xU/3enaZvaZ9tQ2Bb/k9rYDpx2yT
Kyh7Mb3r3HNJ2eu43gfE1pienQvBWj5dPqUtjTDqpvyLAhjyaDDmc44NRJAf2tpk
5DBVc72yfY1RnqOs9Lnla80lqWxWsH4VBK0bbLZXjrEM+nck8fFbUE0cd5LlXnl+
tRgkEU812fBAhfGC21ldV3jkbTKqYHNc4C0+T4P33dX1k00M3zBiCX0wyrVjnEG6
3OGuUhwqF3CIfuprLIkZrqB9IjnzGbkij8Bi+6xRT97kd9RZjjBQf8fOnPG/3NKk
pZuAoQmraqSCMq2Iya4V7s+6rYav1TdO7Rfh1MCn+8hYy7Y8FYFlVBJ5W4/Ok5jP
5Y/eCunGeV+t0OOmsOENEQ7KERald5r/OH4OpQAj+5hz71T47UqjM+WpQCx6GiVq
Aga0ukZMaAie6HIFOsPBGrwyxdSU4vdlNK88D9i9XQBIiOvjec1moenr+ud8/KyT
Gf9tST1Y/EOdjOq9VNuC7Y4NDzfH3ScfTXXEkjm5NTcbEXtsqhgAVugyHDJw98jJ
lv4gAu0y/iCRh9hlQn5H+K4uPWp0GVrCdckQRdTIuNXBm+wYW/ZoiupVaWnScQfg
ivoBiYI+FrfIcC5nognajxKFwK/Mo1P7deXzn84sssbIDFjO8oZCNZff6Rrkpj0T
/VFyVIMp2V5jZYDEkeheBE6nxKsvO4ScSsAB400JwI395IFRVZlqX6IyhanTiddZ
MMQWHKM38r1494hxskfFbcgdTNizVFWQag8To7BdqkKNSAKgjOZJIwQ2tffIW5q4
/ZFUz7uXiOc8gde+tuPIfQ2hxu/vHOGQPTkc1oE+z/wrMAFvOlARoW/t9EU3WxSO
pDugy8qBEdVzIavfjdzb2+SA0+n610Q1AxAasGMflA3r/HxvYYA7+2gBhQNnF6sv
XqTOFNpb2mnL9Z35CFD2O59JTSoAjp1Oi5jzN7QZ0lPfG8ZsEEJgTaYcGvJhGRX9
Bp3/aAAr4pCbNC6Wh7YznLr+qFQ/aH2iMBJxMRJIXIFnQHvDVeL3X/OqdlcQo1C/
ud2QDkHWDuwWRhABzi7Pbu59Vaj0EETMbRnBH0yQQmH5RrHhzG7QJYKR/AcN4w7d
H2wyxpEjIo7rda5ae2UIuoKrGvwQZ2bY6j6vnzeRMK58ZYBlLzShNHelX8F5VZhx
IP31sq5po9XGNfR2HxoHu7HgV41lOjnqPPbgzFqvT5Pss97R7gZTDPui4pglsfh4
ig7rS+wr5XlZsRlkG4diKfHlIt3PGsbuuJbKngZTWup8O0z3MZNziJO7yTuNNq6V
cKba4MWGDcM+bE8N7ITphOrQYfvDH4pGcZ8PdCtR0tRp513KBCmmT1IfKfu2eMZt
bhauNTAfpjyKlyPjCtEQlQF2WtShlXwbtIGX0BZNU7cuA0vDMkH2MlYbaThcnUn8
b8PB3zK68vXBNvLtRwWIYR327zfhqPy5e7mcQ+RrZvhFAW3Cj2p+EOhbPM3sn5S3
kNGDSQbUNYrH/ddMTgkVDFJR5F7rOtJReFzk3iqratbaakvsKpsRFLJtmiQtm5tB
KKecSioh9GqYEwXOqmZyjuERgJVK+hzBqDDsHcYhm7YBd76qafBZRkLqDy0PEeNT
fs+hsv9YL8+RMML0wRAuhQ6ckU6KSNq86jG42gr+A2j/ApLxuw5oLqF/NvHCwwoF
gjemOehacepxGNEr7TEEeva0FOSs+j4gIvENia2dVmcmAjLiO+1m2+OxYxG48MSx
tKnFfroQYD6juXoBoF0Mph1nG1fgHhy44Tnid87rnt3AXi+g1tr5eo3a6PUKHbV0
pFemHLzNRmYiyrGBI7Bv7vMt5zZNHpFKO+91NzbYgxKOyQH1nX5j9Oq9zkvQrSvh
gAIUy2eAjqTz4beG/aOC7Ys/0a2UYcGkkSF2IZjT4/vqOnIA8wQXu5E5bZX/A2+i
MWrA4kYWqohWoh9Oq7/sfMbF0up7PyfqINtQsVShLceXtZcikzFqsxpu1QPIby11
I2oWgqaXhV9ftuN0phAi9ip1fZ3lNG5SeWgCSehwbJxfXFf1RLOmrBcaE9Oimbwt
TP78axiSNanJSVHwduycEzutHQ7Ajav1U0Gf9HpvEm13b11DDuvQe3BmExq7w7Jr
cmoHmDbFATnPJZBSd6614oKcDnDJj3ajqhf0YScHpW448blW3En7oWpXwowmyySs
6iUL2BwRDJdh0vJYnHltd7mG5nF4SozFddddMMm2UtCpPsy8IHQiGFsPKM41Nd7w
QKoft3IQGZEYfCLBre/7GEgoo+i749J5zES0rzttMCm3IAWCg1kqtaqtwrts0mFC
yZwBQdAnLd44KMkh/90PotrAiwiDt8YFMqch5klpELni0ZDfhroP1fanuF9ABCQU
ydlT/gb5nRDkE5b1//jyItWrxwV42H153ySTG0ZRF0abjY2Dn8a6TOzZV6GsoDTl
7aVbUjOjhJ7fM2tQJTjZ182IQZu6NCC7hCY7qC/zPtvbNz8nTamlTL51lzyfYstl
rHJcd/mhovvORB8wVtmNd+eqfyST/8Yoy8DxG05CT5iuQ9p9wGRlDoqUL5V9o1u5
CIDmKL+nZyItwGbuZxoItVRk7UYEbliclwjDFkj4T/glP5N22Hg627P4OYq/Ro9v
Ut5w534qVjYnpKURe26kpK1qSr7tQPow1j3sK8nY/mVU3cYE7PkdXE5KfllTaWxV
t5omLklF8wlDWT5OQUwscegfl6x7SMZKmVhy+FhqPdo1xBL+lsdtZsHSEsuANgmn
LEUmvPEVPmRMEzztUSupVNXUpySqi4fRrRHDEmi5pLz4hsC/xHLRg+8dvVFQYyKJ
lFQ2y69uGJmld6c93cAGX5LnQ8NvrSwd1VQr2gnzYkxQDnjnbLcja/Q8nVlwWUag
kKidwlcJLOV9Un/+3KtGGPE1Wgs5io+0PzXWXTxiiSn5qOdwiNZpQ/Z/Yb+hx5+P
d1hb3vboRewyY2T0H2nJBi4CjYsZGTcerzKSIaLWxAOPLiwNtBPMuHraNVYGfVKt
KWAMQ3l7W9mkDpVTC4beM42U5glSKycJxTBB7StaSEX1KadCo8wCUp6b0PZ2ULAc
8bCPS8ja9h+vV/LBaDKQBh46klHU+QpPiNVUjS5IFoPumkVNDrm2k5yBf6COoMcy
QeAOIKyXDO6ODjnfHhPZz9fvjTmfbFyDsjqDI4v6iEeVknS8ZBdz99vbI8QLhYs4
zDTkud4WQjbfubVBfNhj1YO0oxRAWK7K/qKe3VUe3ZKg5bzvrWWzxfRyqGxZOXXt
EnG2rpn4SW/1cjyy7/djYVlVeSYZ5dULCGvbLIiJGoeu4AXuNvReL5V+C2g9cbk7
SeCK7oeCym/9Uaeur/+CyYQ3bIH6upjN34Zh9hBBiNRQKmKxYl6OL/HGEWSQ6TOc
7G/HTNXJ/hEcP+mN6/sZtwgbbrDOT5igwpDYRD8EtkNVldNh3vg7OD02KmuNbSTV
DsW8W+iwyHC4E0RqT0+gre9tilgCGKZzBLgep5uj8sq+2+2/+CTxmwAAuPtFDMz/
Z6FUZhfddSsNBpR/8SbpTKG12sPVEzWNHW+B37KcSIgQn+nEmYYO0CAzhYCRg/C6
Gs4dedykVN0OXVlzvPA4Y2XkXvDZCHKHiIfcMEqHiN07zB8G7DPCGz2/9bl8ElMH
q4yfpLGhdnneWl6/HF6gekFkx+R9tiFgoESHi2zHW9rMxZ5YyBxLBx8lsza73Uj2
HJ8ELxJ7wEcAr2AEaiWFWVkRCVMYS65dq6biyczRASM26lsaJjujP6tZN17G0ZgP
urjs7IkgtU/2JmMDhbdG9+tS17QmRi7v0zg4Mk3l54ewUC3dua+7hnVOfWDbIb0m
iXCf+DTQjX5ECm48bjq2wfExvRye5FEe4203eBM7VeXY7QDjzBn3vW8u+4u6ttbW
/c+ygtxlHI78mYFqvrCP8F0Cl4STJLfuYZ07/JLDNAGQswza/VqOFy3ANe+YwraP
8WXFaYz3I4emg3ARvjtCO2+49A8pVl/+XIsk+mVi9qsdheJP5d5r1+W41n0KsVK+
X9Raw8sqesURerXoRyoY+oCl9LumEo0ke11y3jkkObm1X/TrN9uRry3Yd+8Apn7F
uNIT9KTa5vRW2snh5ma1AZ5j7R1b4IL9Z445KqY9WHSwJa82rnKQltONFY/KgJrK
BB4wrDSV4DYGLpuCSk4D7bAvvLQjRca6IAWoSaidbKqpFzRPN2i6+X9ukagmWlz1
0egQX31/U8bbUxv6DiIxYMVNlWA5OOoKFPLQ1vtzVD27YuR0Tr0bifMdOAhOdlhO
a4fpXiWwWuxTduCP2Qk2ZzrPfSY8CC9XVxp77CYp+pj44zOeXTnMU0YewB870bWa
WttWKx3r4Sg16l9IXSZZ8x32A44adkHNtn8ELGFpLtwQlwXJtZvchtHm3mc1+G2I
geX9GlcnzubHYOXW/zeaHxxf5Dex9d+9DZWy/J0P/QD3L00t82WivndvHC2nb9Kh
I0QZ9pbohWPBw+jCs1xtj7Qx2fOmviwipKTlJ+G9pH5q9URD9R9Y/jSA85q0R8fb
/Bbtx5POofmQZgslntsecGtjO+2EahSZvDIXBq9bJpDh1DnPTwZcxe2uKMK26B70
PGwaHAK4T1KCVXErn032cl2ai4TKFNtqztHmVe4Oov12tDDAJ/i8CGrXJzLYty8j
9qTN9FWkakRYKpUdMj9v7LGh5LH93vVn6rF1qCB7Vch7gTuHa5q8XIzBCRIEuUG+
xcnvA1HE3rVdBy7wFNZiFI4MEfi7tWIgoZrjCKvlh6F6roY/OfuCCJ0/HgJST6+3
eVTh2m4V75sSENp0RoHAH9RiC+CKijPfjimrCR1Q0lPnwIWNi78s5Uy/w/TCqeTo
U0cLCXUM86BKNMMOmQyz8G0ECVvS8FeA638E6mY8Kr60yDka17WkDy6NcBzZbp7a
ObY327z6wyJ97P80A+gcPLp370+e8FOFhc3WT/fn98XIPK12kXcbOZgi0QqOfYMw
6cc+VHOwoluhAm1g1vS6uc1JcCBknRRS+bf1fxSmyGk1xdckr+TahOmqsg5L33rP
p4u9aMlpOnQ48MkjxbaAJOUX0B/dfK1Iph5z88284lAPf2nydanecdBjScYee0vr
x6FC8sm2PA/7W6BgI3hNNfoPdCRwcWTUmX2Poi/C9avLfDz9NgVnd8I+KwwOAcxp
3QvVHQmdAqhnJKrnd3FyOK6MENDKcjGFLMcCzZ84/QIOcbfUN3j0mSpllwxD6FG+
cgopt4dP1H7vdqne9j2CHSclYz3fmtS9Ow7ecEpeLH1JKvSW9DyOTljl/rqUKCtt
ZfK6eknhTs71GfCdkg4XZGo5typrw7ynCE2YJbIv6SsAbhBiu4wy+Y587s/VtXYT
l5jIKb3c01U/bud6IWD7eE6OJIsG+seEgIvKx98BwyGanLXJikZJGiab+rADmyn+
RrKhAtTrgrgKlmczgyXDfcQhD0c+m6wAf1QIFr+lJvlWlf+P0qpaf01fUwmHXT8A
fCvByy00Fvq84iUyTL0Ax2gYck0fyQI9njHx3mnnJS0Csvyp6FyDPu5k9WqTWzCU
dS47TVPAFCb0mfL25qWwVlfKzXNBuXnkKBij2Apz5leq1CENAoI1LkI4XjYM881K
INySyQ/T7dIlu6thJhkqJXQVB38zw6PsyoeZ9TlyndK93tEQdpuDOIbgsGRWHtr/
ozrtk81WY0SmbOM9IHOyRk2AnSCuO84U3veLJDxMZ5xHZLnrXR4qhFRe/51mw464
X5+wgvl5BMXV3zUFepAReShTbYqxJNfuL8JNr8fxnw64zgy/gqrCtAiBP3MeEM5/
uyxlqMiNyiKcuqKvbQboAxk9Sq++g3VSi7SxAoiioi6HL+wNPa3OKNacdZK2xxuA
xvFNN1+LGmTjRn7E4hEmPn6A5cFGs4pjf6Rkpal+AnVm90sQEZg2Kh+k393UOKLs
ye7+jftuTNXkA4j0RgFH6Y4MhBv5n0Tewv25RFRYCz1KTXU365dAZAtDcK0qXpRC
nHW2v0FFvIIf/80R0Yj8yI3Kp3vdPqXb8qWxhWk0SD8us1DRWA9YuALtXWpT5Sc1
XeVoSrpGrhLTsNpMVinxxeHrwlsnv/tZtVgaRtf5XVmNckR23eDIYQ4A3pBw+aSO
08P0+CU2OTd5F8ezB9fMZr618kaxLO8+urQP/z3jpr96JyJ9sSRxG1LlMDLSpbco
8VArweCIsB1Mp1wrFgL09os8yU9U2LU7MuJA9Fg6MoIGB5wOLOi39Lm553UGmJY3
nOl37VHDqvn4Uvmmjkh6atszkokoNl9byHw7MhwEt39Jd5Y6CpTl6JImX+epw10j
Ou9HibEsUEuGnaXmfq5iIUjSJQkNR60/yEJ3UsM5lmpUCZqkfTaa4Lfs8IFfLvi/
OcpAtlnF6KkAi4w508AI1wZlVJqyQ34Y5tN4JJxv6S25r6fvl2Y0X/V2wDEdfAhl
4yqv4LqFUynBXlMUNShPEcq+8yHv2raSvn2iLcD/N1ZlTb6FGE6CH8icrpcnAuL3
TAU5kaRx0gqhwFrpVHcWfuk4vcqOpW7MgOrdS7LN6vMVp6D2x0XuaxxtrJGXIi38
TSl5nq3aFVaaey9SeeF7Z2jw47VZ8mePp/LtQ06PNdd3WtJiV6YiKPxFqj1KoABH
qUwF3ZfIhFBYTfeIzJ5j3aDBl0o64wDSoXagJrrettev7JAQHrhDOaLcQMD0cjD5
8GOWz/kfzkhGJahOBePCJ1sfXzOnvVvA1JqccUQEngihZq+3wVeQZFCOnz8egHSi
DWnB6VIdnSGqhxzo6xYQCpbdGpkwWa8GS1mYhcQO9GFdgcznyXYAYTXk/27S5937
O8yhdLFYTGxfAvDS7JJjBOGgHpwDcw/mtTjJ7hxVhwZVf/Na13sc1di27wMEEAiV
looo+p4fl9Xq4jWoC8b+ZjvkEAle15NFGQntF4wXA2IdVPqMCLxfw0/m6DsUM/FQ
UjCaSQPoERlK4Scjkkxli77OEjhnddhVrN/rNg+L8SmqgPp+XpYb573bwTH5/Cak
ic9sxGg3XbQnyJyGaUtUg8UMwEfAkvgguDHpkJf2VfSxtZmttWiKgGfeMl8oBm9D
9dbH3rMu+35VVt+2PcCtK60isO8g8a+Y81z3a/hhYW0O4VQt1Jrx893klsIyCNUb
s3JUF+YvCcx2SbLAXqCZmkaju38r/9dQsaPeHj60yZ58mQ9kON2T4T3TazcOa4dU
Epmn27FT8/G6Td4CnF8J+865SITg+4WwUUtxr0HW0gLmZwqYvoa0cNxkv83fxz3d
MwJvG/UTYLeSx55UMHksc4m5/QNR0CNCA+7pIni7ZkLqbPg4UpkzLQa6BrV31FnY
7BZ8EP43E1/Lkmeyi2yGZp85f+fzZyhXLvvD/dNNMhdGQsqeGiv47SDXIp0WS9Yf
TBpmJBUB2eyR9zTM8L6QDjun80K4xCbjvMsigCes3+2zvEv9Mg8HDr6Hw6B0eF9Y
wPdOjw5DpsQA3ivXW6JZtmPA/V+psMOLBF1PhKyZC1IUHLuxZEiq7dY9fFGcw3D+
MozKkTl5scn58Hg5Lku++goIgQpm3CG+kdR8HshaCDwYX9r2h70GYfLN1FpF6eRp
9ur+kxEeDp9SsP8gfeabjZdEM50/v68aUF9UuUU9gOgqZgVENSJSbuMlMCE41N+W
hEcVyNdKKd8eTMPjFhX8o68yYrojbrDxR/H1Wmu3ktl2jmrhGL0VCD7vZR8BlaEb
QWhQSpjnL7QiZ6ZNNRW/WOtRdi7b4PYWRGW0mVABPztGwqin0l0Sghovby47sO+f
6U1tKnlEdtI0W/rNE34adzRjNGxTXgwaXarHEInwV30ZehJjTGa1VxBwoxsudrZS
5ZFbKsDwdQZiifC6DA3PYZwINfZEP/asUFhabhMe2X8FKU3l3bxiszMcL07fFNfJ
o/jhEF2W37gtffucQnf/TCONK0eyg1C6ldp4SOQIYOJNRZp9Jgvj82r7fvdWyIe5
vEAi65DnAiJU0VUEovTQpTTKL76bykO1iTY8eJq8JnIzD8htSTW2l5f8dQH300Xg
MoCbaV9HszfVnTaApVxevVg6yktbNk3JGQ9M4dMHrMU54L6pNxRRDyLqPUr3jZj8
3atl1EJcEerqnNbJzAeCpxnkKWnrAiiCHKO3SEPytdX+KAb8T/AT71QQHmIyQJYR
y8O7RGD1oY/bGEHsihW+OaN9/THgbWPb121CkEQTIEP1GNZKgJVignsfd5PPuQBR
pint2hy6o5fkEf766bCcFV34z/FnvNap9doq6/FrZFhGJuxznrQSujBPd1z+z+Ih
lby+uEbA40zEwPSDAGik7eTD6QhcXOZLMajuUksEWyWH/E9ZjHKW+Kbyl9UvNYfP
wyF69ie7kjgKKYW6jmy0Rml7LLcqezJt3HbSNXX3Anxym18TILQnQw1yO3+SsX3L
U26T69fdgrvWMpoUUDWxDjw8kSkJDO+ALt8kVwgOXYXtcS8OkFSan7w7aHQium8U
jvGLp4G+AsPuacHgSEGs+/Sy8LxHeI+1FzUWc2hX/TLozfuIsFBaOk2HE8IQ0/LS
hb55hSwiX4CjMpIHGuwnDwhucN4io1ErMb5YusJn8in4jAJx1Tj40Fi1tChcROU5
jYUR1FynQXsx7P1brcFaeEI2DFagNRmyDY4nJ8BTK6OjsGTHAdKpaLQohVZG2Rz4
6JIsBwMRU2yKSmYcxAzh+aA4Lyo9qK0TloBSPoD28iooGG2f3Xi9SQD7NOFOCuse
Roa7x1KxcBuDtDlsWgEt3qzaQiN4Ta2EUc+XIqfNOS3GbX/b0Z+hL90a4+qtounI
lGJwufZvt6oIUBB4nQlGwCV3Fb6NvWzNMxMinNXLIPgGjIRLoehfFlmzOkN6AUmm
GY3U3dOc2TWA+XgDitkLEYX+tFVML9tX862agOJ2ev1EahM3+ZTITre8DAWJDUwK
koNI+3YTjZ/ZOcvx898lh9nM6SiZ49tdwQEq5LTGjJQI8fP1mRF1nCtfcGZXfiEg
IqUbBjuJZCXqmx2KDPJLyd9LYTGRvoKtFIcE1ZV2YjsPL++2DE7g6JlnMs7mvtRp
/HNbtiMaZ3Fgl0NDpCAaDRPL74XCil3z+xZbrEombZA6JF1eDzP86Mk3I9HpAbHF
EW+DP4OhHzbN3fhlpe08OuDjtaf6T6MvzfrJcKTfnvukQz+HNkiuIhM1mpZQ/B1M
UxNApPkVUExgo99v+wWyn+3Nx7YUXH4LrLzMVNQjSAlIwE7wQEgKI4IfDFF8kN90
uoGkti/Y4MwZeEtBbmysshdaLJQRLiuRXqJhwytgu1vg3+JhIz5l1m3W/tu25cVQ
3mRRzJ8D7Q87DwnFORChE8p3tXw+E5SLmDilAW0qBHhMFQ1h3o2POdWnP3gibdCd
cRpq1WvtFNWI+VEa5jC42xyZf32V/0FXldT3Ot8tUCybnTCwV285aZbdss1iCToB
OAPkWbYeKT9FSw9Rq2sJ2bd1Xda2G8+Uudm2pPtXETeKbuBhyEbNcShz/UPyZu/k
gR9Kc7n9xpmav+hIUJvdPTxjKCM5OPb7m4LVRlptfza3yFxgMFk3JSl1TjNpotEx
qmSYU/9TmK/VRvz9NrqqIVQwh+WI3JD2hhTVAlA22du/Cw6YwQ3NiwoovI/1ktBH
+Q4vUJycPLhF+0OrQxmDNAuMC4mewVq1GMWRDHgck+iVbiz/qNDM8Env5FJAvMQD
GfVCLMsKAQd3A7YCdAfFJT3sVvAgUQpDnsyOkLxttAzz6f5+m5ntcxVwueSYsHmU
7f/WoF6E4Dr6j8QSPyzgL2kAdFLd8xvfk15ThhFePji4HBLREF41T/jn20MgQKH4
yMFX/bHc1FHhPxtLZVem/Os6sJWw18VNP0ezOQfcEQiVAFpTJs+wuq53GALBigDV
RT9lJa6iar+h56xnFo0TgsEcUWV/iF/cjvMsQKQonqusGY/Pl23xam95cBUHHrPa
Sf1eDmnxljx56s7dItr7/7DFoPPXqYi+9Hwx7iV0OpIh8efROAUEKUYUiVscg9B3
qEMOwdbnJVLUQvOA9AhayurlO65DhBrShVHESOeK0G0P5bxbGee/ZdiJQLAksxkW
2aF0rrGUFE0PohG5kzqM9bUnuNFzCKKvhj8r9N76d3Gq5ngCpSip9L3WittUlAda
k8THwxmn3rKVBzX7zml9osTSHV7gXWKDDElDJWlIMgI8LNHlmLIXClqlGXFy2z66
H85/As8L4F+geKP7BLSTtEdufO6bTzD+6NhPkEvDOCAhqzznQCvW+6SVLRMkU2hS
DnS1hDP+BnSnkP2Z/Qgdmze1SCwIi1u+BMK52IHc1M+CZi9XY1gm6XHNJwn2xh+U
hH7uc70oisit/nRd/Rk8fjvHHknL3z4tNKp0SgSO80L/3Lc0W3cJAKi4abqEHNI1
MaooCIocBwXWw0UzcQDH7AY8Rpeg0I/H3fxWem40kEGrbMqMrWJTTM36ja26dzBr
n43BgaLXID4zb1z32nDIE1a88nxABFTuX3DPQHxrIc9I7omez+qEBo5pKBlpk3kV
kEyHdF9201kIxhL3ucQwWeTxO9Vwa9Aku9UNVR/HUDd6vAZc1ZotV+bSjJg8k49O
b0mrCKVTiXW/JXGlSs/nHgAToYjATFj5MF5TUQs8HuJ68p+dXq/JpVAAOgBJqgA7
LSRSrPmPVR1jnR/RTs+Lv8AnNJUeE0cHQmya4m6AtoZUPiPWq9uGthtfI/V0cijx
UuADUOOcfxmoM2vndwWfv8JBHrbohoF31gnpB+Cw+DmQ/gEk3T9poGKnbtE1nC44
D7PrkmzIR1CsSWyXpMxYs7vLclZOuVWh+cOJ1wd9iNBxaspFxbq5OeOUTNDlpBZx
cbECVvTRhSMh9YEtHTorSQkRnHNZ2mFxoFtpiX9BgpttLUSHCVLRIsJ/Ujw5w2tk
BqeI2yBPjiwqGW3G7cSnPuMC/WXBMmJc+zdpucCUKmp4YMzTEHMPUFuY94RE378U
D4gsZ0SFUhuQTvUU9iaUygOkDEVjrsI1BB+Cxve7lUnFL02ZLzNLvrYA7vhi4OHb
IKSm38AIQLxAhEzLm3Att803u03PlnbmMv/kBnLE7q1MIexUOMpMLV+b5YyV+usA
R3r66OdzOIcfoWaxirHKYkdty/uVwu6TrbF0u4hk/oNVmNj6hEsjpZRjuvh0fy4z
okQKcc1mg2Hlc82jkt2y0mn+hceVDjJjXPVuesSL+Iqv5ywMfr5faVTT8TfZM5rZ
0hX5z+lPHxJt58vpoUZQxt/NejfPKoBj5QWXGJ2t6Fy7/bgjpkct8NVLSDfoO9mC
WfKAdIg1f5+kXtSvnAYtyc1ZVVLS1jqn2utHRTfVkSru+oWuCrSmDebCzQhDyAag
SQitkZWY8r4KgxD/F/pMoM8zILCCFWTiZ15DnQjJZGRRLCETdM2w2Zk8gj/18gs6
N/cesByQhdWckcf0pAmFN0HfUQdhTK8uNM7Gx+lJZpIlML3U9zFz/ytu9uXVp/0p
PCX4U6G2cHnBA3yUvaqAw/rJza8FNAigNGMtBHhquoQHcNFtkgMRrCVeTuU2KDBl
DaKjdGDzQEycZq9TvWR/DYqV0/XejBprqbxf50AerT4gVGgCvioWqmDCcnc2IqVR
n/g59swi4VYoSI0y/92+2xvEoynefaBcQexRHW+BONzOg33d2FG9WnVGxBD4Yl5w
+vHITCNuycocQgcKTGPoaBUJMFmxKkvYbJUNNsyS6njPgdh8kehXFoe/g7SsNzku
4WUyeqAAA3fZWRx1x9YF4Prrz5C8T+qZqPJm/VpYmp34sqpTdT9CmxINswpuHGVq
k5GLB4zXsrMzI0sAh7euNw97TTO4eKOa7aadD53XZc4ibe0op7GA71KmY822T5Na
fXnZjKrDnZYZ5/HYxR5YJ28Ta4D0Vfmd8DKybKO4ahlA12uoj8Wpw1pWJgzfYXiM
NO9uNkO6Zjc7j4OnQet9wozGzirIpgsAbuboCajdyKR1f5ZiJKWGMKeHoNaQXgOI
UlP5d5sjwIJJXHIIKOiWeQfjIVpYmVGiSlIpe84fcvs9eAbEt/Pqh6qUH0sIosZO
ER/pq0FqjB8ZYdEYkRVLOiDoCfYW/NMgW5lC4OEH+SxDRBFIxRoPqzbxm/FN8nnI
LwGFUXz+X544koL/HsnF8XiaqfLxDpluxsGII56pAY+LUSvMlZ4luRK8m1pjUMRP
YNaqDGPXAvk+FEmg98La4ugSND4gNXgPghpbv1YadceHSNGTYc2pe45F2j3R5+zw
KcgdV417AGjBoB4ZdZvYoUGZgW6Ftntk4Ixzfho+8cX6OpRy04HIIdVIqWIK7DQi
vqZDAzhpB7F8IadzfW4VY4dHfQG6E8jj3sWGm7E6P06/gqK3BRcXowocMOjMTtfK
xeJSeG+Vt6qJ2Akpnt4CCDAOr7MK8XS7nRg/UtCawHtl0p6uHyl5NWrVSeFfewzP
cHN4eoivDykrIy8JFw5OKW5GVwvpAT8pfr2sY218DjEGuCyde4QCpX4Cp8lX8wh/
Ua+ePxe8fVXo6gWlt/NfDHbV6RBgLFQMFlD3TRUYoLqhBFrnv64Zm+ihaNlHrjJ5
WZ/dNRR/rOvPjCo/Uy9CX2sldAVYFY1nYQsiyl9NCMDLIEykAnw/CBtX8d2YG2NR
EjD0qpyo/v25RcWjVV6pXDQIJYGFmIvWVERvHg2EHF2uJjDUiHa//kQtdJwX7AtP
XI4NH6kTMwxMn2iYwehMGwDrxkG53muT0/AZ94hoUzTiBcj6nH4fB2dvM7Wr8XG2
GWKKD8bvygiyoyKFQPJzdaW5Vk9S/5ZbJ4FXhAgx8HDp7BUYRISTsi0xRvb6EvXz
3hgr/GpRJnKRKLRw3MAtc50SuoGOFi0W/q5s9aWnAw/Bz0IH1SiXWkgytSEICQOK
+7APNT9yrpvEnQY3M2PjG0Tzn/TgLXFZLVaH6obYIGQPTs/X1lS+inaYg2TziQrp
6Z+L8JpxM1QTFfesYA6g2NCWENOriAdbLKAWzHUz1Ig7C41MmStyHGEQdk9l8euZ
8lUzLryMLZoCZCzGeiDvvLGjalLVBPCgGCv1b3Qyz29KZSMk8odejBFU8G6fJWv6
adW2icZQC1YhmeJ2rX1TuziihR7UtQAlRsccJDjunXXukwfGaXqqCnqxnBw9D6Mf
++Yx6UU1uspZwzKwvHcts1RYqPbALQmfjrN7IlxHvO8BV04HtsU0JQqdNYdrXCZF
kodM6gaqKBTtxo8rOoxi5wWpkDeSmzIByOhD+qvkk5a8LfwpjxS6o5+FbgPtj42m
doKN2MDFalv07EBYkS8elJMVDUfFLUobF05f8iWGZm0pp2aSiUbUnCbvXpRSm6oc
SAtbFO/87mea0hPyq3bIEqcXz7K4E3RXvaUMQ3QNv1wG5YtHiNfQ02mHCPFX+Z9P
XXxMI1dK0dDwqEaJYKv/1IIU+EMK4YMw+UmG0tdhQfvAeco9aKRqd9VbqpMI1PIU
8od8Zk0se/644mMFFKjjmjQ7/9AH8BliqCY1HaK0kM929tu2eeGChsBTRV1DtFop
qD5FDzo1jkUBawR3TxBfFuLx2PJIV6FYUhzpssaU/gOY+ZscfhpxN9zIMBPOB+7Y
slYZv2xYBk1jVA1R2VTCDymOEsfAhJD/ngHJ+fcNeDwbOjpzGT4Zn+nUcuqZS2Y5
zp2HvfmrmmDyhDaT3RWUg4gUqAtC45zCe57knbbApsb4KfvX7NYGGUIHBpXjiWp5
UYe5UuHdxAc4MZsAqM3JpVFqmxeVSae4Z7q31FNAAwSt4ljVq4xF7DKFsVwS4UdH
s+iGxUXTR1ddjHye8iS/V19YduZBqObgeB78zVWKPuhgIi+9HkbOa9GAY8HxDEUA
ZnKCFHWrMRhs6G7fAmTCLdEV/bdH+5meFoYCWK1aKCeqOph0JqciHlwsHw5JK3PF
QqXE4lBBplaswLcvzKLVcFFtW+utvvyiQcOsUJlUGgH7SGilB0WnQ5Bqb/nx3yB0
kYTMI1IvGHtdtPCpDdFPfkagR5cZDcKHnw12nAv5dTXFK/gvR0OgiikAUkjm0mzd
3TGDOWkSyZ+kNOAj4mMGxvBWC8PN23xNLSQ7BDxm0gMSDMfPJjd6Hxw9E2vije/0
ex4Buqk5Xn07ZaRc9JDYDnFbHZJ7cVoHO7LiiZrQh6vMigsnsZp0aPO8Dpt2Jzlk
2468VhQm9Us4ysg27qji1Ys85U4lzQ1bn59H/iNu0t1sIqOxysHERNJ7yul7Dk4j
Jws1JS+3Sa96KCpyKOoZcRvvkksRsDp9G9GVlFobMMia2DTDG7dSLaqzajcHnxsW
1CZ4ZaqikAcOnZW9vF2thh4/G1p5e9eYlztO2mX2/gpGPPy4ETPujLoxuCzX2SWW
wQ4LhoyWW0WeWKXNo8SoWpxmBosLESxfEf8FTAP3RHBh3XoXdIoj2vQqWPUO/yFy
qHMS68uFID/wQh8GnJIQ0HoIHZEzGppx7tAx5r8RMmek3O1YgaTZ8ec1lbq9EkOV
NuCCzSzL+AVYAoyoYmFMu990KIujavnCAg1SwFUECrXA8ZyplNNyBYzGQ1N8DB6T
Sgnju8IOjFNgiXuZ5SNrbrUMLpNHIrFnQGWqj2luPeyygSGpfYBnd99HXsQTuahk
LJIDC51B5sFCh5pJg1ZJHw/o5q0+TuJyfZKytJnb1oj5i4GsJHoHJJ5VPzY18ILv
TQ4HmMx012XyjLtcXzlTuKu5YJHzFNOdAGKbn8x0aggZ1juNPnvmjIDqmIVj+yO/
aMWiImbeovwaWxHJpI4TRmcd62A/JFjtpEodqR8+ma+0Qg6CNQ/5FgEDjlsKkgjV
Utuo4dnssnATMoGkd0I1lNiMUMLS5rSu2kq3bA6s+Y57g9s0TmPx68FfnqZOj9j6
88FI2odjZnFkGnVjw5DS/YExE0X+t6p2sDYklGsjVQLfiBFvXJdHBjNQFz+2Szmw
r+dQ28NdY/rsa11lEOSMkA2xR1AL+AczYOMcjtpaP+WhWh5EKb+V0roivP9wSc3J
WuNK2Hd7L3zZAqnw6ft/2bWrp/jWcZ+Dj+eXifNdR6Kpaj72d5zEC13KXn0pVsdN
wKeENP4ZrthtDfyAX0XQElbGAdo/A9U0EX7s8L2WMxbJGA4gP2qeEFiFhOOQvHzr
nx17cI21dZWnP6T8x/Dchr+YnSgCw9Wgs6zdPM86sHCynp0atyO/CZaTEdOR1CBr
y+BFu+uxY22GpBzQPRWaefe5Io2dTCKGspeKLg9ACRcTg7AkfjR60nSw1nuG3dHW
p9zZsVUTCL+NwjEo/qMSe7HXLExNOR558ChooQt90EfwzJzqSfXQEKj5IkXdmds/
lrOrQzyTRUb2SgC/8Zzuhl7XD1WG2neMYCkCokrfPT+BB99T4WxgJyK0uFUPrck7
FPHr/A/LSL2CVmf75+18K+AWzG9+H6lL7S+/mTfoBBb6HGcIIyug419OjWRnElAC
G10NuBA2VFopjrRX+nosQuyz3c0if18/ohd0p51eesqRrWuPib+TTx5GWIf8i/OV
8T1xTsN/1gfA3ArpeIA6ATKWzaCmVVaLz4E2LVJ3Ft9Mc8c3ZO99nbiq/0gKUZJI
/t1kb/umsA9xc2W8nMHSOEHpahWVqgCLWaa9gsjm3YphnJjVKdl94yN8CG1F6h3i
zFvPQY+RDTdYeiejxyWYblaISIrVuupcCgfx0y+aPmeh48n08SePxH3YkG8dCQLP
fULwUT0IwMdjioTU1k/of/HYoNOaWETmQz2GjKGRa3+QcDLqix2oFYrrhuIR+01j
XTbw+BQNq4gqNsdqrCPY/mQGkkMXeIdrqWG4p2QbUl8irg7VBOnJ9BgzTCHwfts9
/IcjVDOwxkcQf5bXE9YT0jzl5dgApg7WFQLasngfns2Mhmvl/1BQi/ZbktgPDcjm
pGwNIWWp+Ce5NO6ZSmYqCI89KRf+YcUf5tb2Y2Iof1EOEn2jKPrA1mZ99Z5XLFEB
gOB4LTitK/4HpVHloz8DNQ922V/HmM8X3dWpKh4HAUBIxySZ/xAm8iWFRI8r6tF7
X9om6SoqaIN5qgfnJ+p2Ls+ZhSe/Y9HWSwbOGZm+EpSZqaBAQJX2U7cWWDUcgjWE
0nIzjXXNrI3Bd0ct+GfbjZYuMPfVStqC08nbAQhmNQy0CjYj1vNuV2psxtUy4eoO
Fcth5rCQ326tqSaDOZMSs6cVhRVfek1X9Z7PHE6hqG2oGzQDDNCWii7cjed5u8Ym
AMwJAhAPWTLV8sF1wVuQLNfJoVFDgXeTEg2ROPjQJ/HJWoaJ443/xXlyyWmKq0/I
azIQv6MaY/sYDMLRHT2PuS7hp59TlVYGnWwtaLja+JEi+llkuwZdhInetIGEUjPp
0X8z269QA7GI80KsDLwqDkSFiVwPMpYucM+b5x5Pd2sNfk9yq8xBc61R1r+F3KX/
GXsDKdPIg4g7CfIrkBF7Cr3GTxy/TcVriGI+u9wfxQLCJfOXGl0kKXA64C6NXvsJ
LcaBJIcU0Nee8i+fKm2FwraGrI2M3EYFJsQ5ZMgeqIMiFDMlvvV/LxkWXRXjYrT0
5VSJEipuTapkK4iXBIrlors92jiqgZiVrPjIgZDZoLa2yWRf4MNp9eLBKKreyexz
H671+iRFrSVfvpVYxNuNT4IqALiO+JCAckICH86qC5BAXJO1hYrUoJnSDSVlGA57
D3bedhSEYf75AAZTnWHu7dL5Tz8gkLFUxNnU1Hb4xuZiIbVK3s0tq4/4eiOmeuh1
1dMthT6Ah5ZhBOj6irePusu6or2aPZzSKEmgYHB0fHAMgIcZgKZlCH0lL1vvzPMN
impy7ssGWvJrzGI85B4GHaSsk2xDY8ATmB3MFhfvmyxNnXUIK9YEiWV8tc0OvmrV
mgoojEdPAYh7jxLzjnKDcTYIeAjAAQyi6tPcnWzXPHeJWxFRg9eLbz3YnPQ2+0sU
1zhhyvj978xQdBdFFkQ3Tt1XsaY9SFDglxYHexi0LNbFkoCQa+2cUqZPfHwMUhGI
oGPdn9RRa+SQR6YjzpxNaDe9cWA989eYQNV53caegguoCNDNZbLekwxEAKBePu12
yXrTAY0ZcBOBWrYzfBMtjxPv95V/7XKhW9ULIKGSMuIUgr5Uzs7JXSHEo98/iJNK
FHkpgN/84obsi0LvctUAzCSM6ELu7JdkF7jq4prOuHOmMPK3L+PK4faDQS77fjrs
qvv6EXhUegEMfoAiVY42k+dkZVQx7pGUQ4+9JGr+edqR7oVC/yFRNtT3olfRjufw
TpddMtXGWxaw8jqRDQxMG9uYa3LmYvt+cStJWnELDOOnzdPgRbpabV77QKJVeUiN
ZAh7dxligpokSpvVoqS727oUG4B/vNo+Lg8gnQIf8Y+9Lc2sS5vclG9I+RVWMvJD
d/z9XEylK2F9A0Bi0Rin4xEPd8BzY8uUPkpScIB8lS5/k39u7tsC4W0ZNe/ALJ6F
bInQlMTZtXghJQ6MiUcEqBc+20jv5msLvSKU1mLnFl2oTHii39CVcnXqKQVJLk2E
PLy66h/tz83z+K9h1ITQbtOD7wKFLCHf2JnBix2C/GaQh22Sp9hsK62HxRCV01Dj
nCDuoKQ6ATJTd7jkSgldNHhU9H2x6EI22rIOjdriGfyXGKmhzpKDX407mJk6Keuy
9WQFqTD3g5iLhU+jUd4Rz66TucQPaU19XgdXVj3D+Tm1YlgX3S81UTsTBmxazyxk
Q240FqZ3VlB6wTJW9cw0RjDMpraVSkHZquKFgKuedNlXMNCwztPC3ZuSRyAWiIll
xBAWufrdZACaAHdCBWP+gO909eafOg762gRKRc6oGwwbQduMlF+YfR4sMRg35Bwy
sRW9/QTCBB0wFK/q2DqsR7acsEZUINrsB7oYI3ifxOyQLyhLTzxxUQDvqdSacO52
eSATMNuyXkwYI0ks7oRupsnm4/rxItgONElW+en9yPsTSpjux/QOheGtMGTHjTU4
356x4bmBkUxmpQnHKZP1Blt718Vq6JTVL/zTYoGJx7vECBqqIjSLKvGaHKmSkTe5
mVBmc/S8FrmT0RE/e9MI5r8EzEJ+Tmheh3580ae1PFqHYa/a5HMGSePFhadDehgr
62Wg1/tT5Ceo22lKT//FHk0tOiEdKpYpd5PwHH36UDBt8jw1sJB6MHU9+DjAXTfi
pSz4oHpwYfXKwmIXkV6cNoZTFAiY9WQcr4wHohQcb7PF4EhKQbis1a0tWWFUn/7A
lvYXnuzeFMh0cWf3ReFz+SNBXttYGSKYhUTZD6HJnLbfl7MrXjFjM1k9dheOXVe+
UysNMP9vWJzx/sElNdLifUEoLBLpj0wD4M87VkV6EaelWCqZVSwT7dm/80rCDs+G
AoJXFADxJ/q2aKvnOIyF1ZwH3ndvRDQFs6sRqmArQopbVj0LBJ30aM/k9MXA2evw
PGjuwNIgnnwoVif5qEzYFsBUYyT/h+qr7A35mwqG9HBwiAZoxeBXOjozSBhVRyYU
WptGA1QRq2P7zuGoFt0HuofIdX+mwpg21beSflU95Zybn4HTBP1gXa3yoLUn+hMO
FBmRL1gnk7Qq8PstalTTyu4KCzFgBSgqC9gvStqzbMq0/OHnzQ7A0A0tJ7NDT24X
JF23v5cJCbzvWg7ndBICDdbZr9xia+53gNAaYat+nrIfxC4o1rZZV+gFtMokxtbO
aZe0DJOCqVuyR6peDMamfNiximMmwaiuaIL9S188yeUF7+eiCZoMY5pT6tbsqws1
415FrtEe+26gKdot06KTVNWS27uas/E1JJnvv2pbxQImvHR4jxFypzuNvQsEeEKB
mTIn3vXqBZ0n2is4InxTOf/Xx1t6V2bsCEVMJpKuhvgdMBojKPaF8NwnCmdXIvmc
cgs4T+Lhypa3YALh9F2neA3oRNPgJqgW5DsDpBaXfZ+A+XLHmT1cVkJrqEARz6zD
nYYLp0JtoRcThATbVFyBJ4jS0qJ0vorkyccbAg+dfRqJN//YTfXiFPAkJMPUnHf1
t/WlKAIMHGRzYo3LTFj312YBt0qeTyfR0OcPj7Tx+e1IGX+yR2tvxjrN0M1Pq/ak
fFIFDSmDlj2cHmXrXlbAHVpYqVy6nz/HS6HiEr0Hpb+TGZjsV0JznKrri4k56D9x
z00BV16pP3mPK0SUWnm8y59IK+MIh5UAJEcxhvrZ7GhtsN/DKoU4D+NNMj3EL1ln
OMStFhjhWHCbva2/2mFkFyKi6ReHQ8SXsQvET5Pl9/w5bsVXRKujVYfSAagyH+gi
A63vKRrXj8wTpJtilzB7d1u2dwaidYprXC1elCSsrXGocDF4DK2lRgkL4VldRUB+
rQpAOIaPykQM+GhH3SoL9QsY0bpbJOVV4AORYxByvMw3nIiw6F7o7HAiCY1eZil2
8aEUh6VL/XrXwT0DOtvD1Q/Tx7lxeeMrrTgQx2D6OGMpjo5/c82fx1Qjh5p5ih2i
Gjht/rhB9DFdBhX7AOPIxSLjqaq/XVzJBVwBwpKVUH0VdAvBnMoNeEoSG79HIsUq
0eJoMxZssIRrgY5Q6Ijs6VmUnKuOUySMtK5q/bIjtWluISM5mGmV9RKSC8Fmv9J2
Ui4wtjUgBuomvcHogzVWZ1+HjC18w5/IKpZvxKJsFRNEOUPVjC2Xcg/jMCzUfEoq
xO6swtoyLoJH8eJ7R2so9vin0uRrc2/9KR1kxJI1likioBq4qNjWPCfHjHUIBK1V
loFbh574CiLVoRwpAh5kMaUFFJNGZ0rW2WnDXKgz79UybLigEuN//MbsnagpAT+0
4HKyFCr095BakMvHs7m6ZprB6hr10ZClHmoTCjADwxvqYElUu0kVo52Y8OPWwdwG
IytdPT+gTlPVcdcqSDKXwEv6I+Wco6oOtwW5FfdLGnXLaJZclmKWcWcN0ZCyjOBB
T+ZuYdzR4zzXXurJRHvnI+BSrqquG8KF+fWe9t89VjTHYliFZaUCDLjZmT7VI62A
LwdOVnB7u5SPB44clp//AEJq2Rak9otfjAuOwr2A6uQzHt92mHRP11rX701DlNlc
ie3aAhFs8t9piAYpABe0ubHwMj79YcVi5aFgjM511LQqBu9NtESbTuEROVgHpmD7
z5lfXMMy0nP9I2zOPSmCzUieN02OlfV+DXEsE2YW7mwezN3X2zOXsnNGohMpJeoB
cvbcFvU+fiorKnvgS7biqxoT5toxrKdyxRRq4CtBf4zfk3ponJwctITmiZOZmhw5
1XkDIeFCEwA2bqY5CipUs8sk9mvQjPPs8IrFzapmVwTLsWMnkpN1jr4ajAJOqlha
T2X4/ErAYX1Dg+3jFcghj1jUuSo+D7h9B0dkiAwQwpZP0e/pgUfvP8vkAmuHh9QA
7S1luQC85ZwrxtULxQAsjixcWwe7KAUyJfaHmbzmPvAhgdB3MG2Hg8U7+yKT1LE5
XqFawW+NdhiFS7Uz313nJTRC2vNuZAp5dWYGfk8o8BpzpHtWgaCHnbGm2AnyjnEo
Aojc7/kz6z7HN8R7z53T+qPIG+jKq9t29Nu7vXwVO7OBL8El+n6/U92KdYWhLlSj
pnqkjwtYNjlQQTbVi+0WHc7wfCztXaL1Hb2CpPVBLL74gz0a72VFwKZOiwEsnbRF
hWChdMhfUEfzfaW0vlY5psuGTaV71x+Dt1oQKR2tZhJp++Fuo9M6xKn0DpPvWnLo
mQ1NkfoWi5USJq7tPY0rTe7xSIdWHE3WdSAYYQOmh5zcL5uzykLtmH1MjvOcqkpz
s8OoJ43vaUzOna00jm2ydqj934005tNO4B12Js6oABSZgJKjhJtkMHArg14vBESe
fVzlzHCQrLe5ixXVpJh2SvJNu+jX0gYJI/MOP60MnJcpVuTjeuslU+dQVrLJ7ot1
4/Sbdn2Oecnz/KXUtztB9RbjbTabavT2sHvXNfIpaLvt4pIJbmVzzuTTCGlHB3MK
NMFtlBDXdYjVXHNW7ujMNfhS9KSSD0J4uUhzDI9tFZDjDwvYmbMyZ8GJ39ybCQRm
5Oa5qZ60GR/wYkVZ1mtNyciK2C7QeUuNRcVKs5uqi5VCL/Wc8yveMy8Zhd77+Sgp
BZV5xU9UcZyW2If4njYlmbq3ltcf7lgo5vQoC3oEArG+6HTsP/hsJTRflp4bo0Oa
bdNdDtORsK0tlSj0bwl1TTS8z9OCVr0nuBpNeKurEbNnJ2RqqM60lPYvzKovR02F
PlU1hUHfod6b+UfNkccnbGQK0CFisT1yAKj+wkX0MtYkd9PU8QuaPAqHQihH3Og7
p2/RhUQSNwTGOknRrqqont7P2rnnQcqFYF6CI+bQ/v90GAYEbcH6P7GOnuNyJg1q
+W2huoZYlvnSyHyUIcf00TKmUBlQnHewJogNDp5YOapxwv4ljU6OYX1gg65x17Bt
9u6YdQdVCRtVuWQsLvM0eZRoayJInS5hC7RlBpF53grKsxBL3M9eGCpVdd2dg76e
qoVhQNZRBO0+wV2VekX91xDKE3FAgEB/h3diMdpTEF9BQxaQ9ngWcFkslfbffosb
X95ZRJk0O4TSdXqOczvnsHGPhCcy5ldje0nkeoorYBKxJ5KtPwOF99LouiI0UUUI
vDAyh5ZkwbUZ2e/K6pFMfaboPXbm0/gdKa0b2Z7J8bO++nfPDETLGJOYeklZKTPA
8QxuOFfG61c2Fo5ZzkWdkj5mW3zfDLf2oB/3Jdm7I9Ln0Zyz7XwrEk4AqhIgjE3w
14e1VMwFSiN4WSIjPegrLSRlzTxBXkPOZNlRaBi6Lo+YTLmeSpnBYCdgesvy2PjB
zfUjeINc1ioD3iOcYzRUY0Rkd4pzi2kckeGANCMjC4jOLSgmjxxe7mTMGiXHxvq2
+f4kh6hRx8UAR1stUw7v8LaSfyM0iK48GDfbVAORT7H4KZDRGCBPqtGF1cMYFsUq
p6Q2Fl5TXrZLXZVFuaxGTaISEVyhjKqDX/sEjx+4Q+PogyVmg9qnzvgtct+6pGk7
h9FDHx6oqccMnZxCb/IIl54ZUMqANd0MA/2TUtPu+BjEHXq7kv3Lx5QZf5yU4RVR
cj27tOgJEdn1ShrXycBy5EKKgoHGTfUEZRfBLGYhwViwHOawOQzd6hIR8X/4fA9f
cVKRLRRhm6DR4U2x1vf1gFf+C+Gd01aLSZeRyQB+OxuwLAxFwvUfZetzvGuDa6xQ
SPkFTcWoD55K7UeFy+v082zWt+o8ctGrvVO3DzLqha9CtLOFjw+1NlBPEuqzGAUT
NF/1rMRJXL9vJ3yQ6r8gxzqCz046znrPVWBo/mgAsaGCqLems0Q6Tau00G+QD1Ik
wnwZKNAIiuuRzxO4E/Rgh3MauFB5Y64T0SfTzLfjAoaUYCJ7NYHLNip+Qwe3lDBS
GdTqb7mwadkXtKVUZul5tdeGrqFAjzm+4vk2otMUmwZwpoVSw7tA3RQESZZlqDcu
/Bc94ePWzrYf6XSWm9R0obYeynlZ2BQVZVI8X6nuTPoJzhlX1bV6ZrfvyMQUiJKi
hD2o8dwcazcX3BX9vuyOCQobOw3tL0daJXL8Ta4PAEysmZtQqJc3JMgLwZI/utJ9
pOGNd74RE5HLbx1MLf4h6xjIf3rj7LFa/znAvtpRePK10mXdNLbkm/kNXfTjtLEX
7pZbUJR8M8u3AW15l4WqB8ksY8k36EUrobHOIdbmGnkq55gU1A9vdleBFsDBgU+Y
YimxiJYSCSm6AIaABkTA33AiZ4/9FMRmEi8R16vM84NxkGkKiajH1DSarXf9aaNr
MTwR2sG0nIGBYNyI7CaDPcfs9CyQjbCu72ZVOSlk/A/vViDmyVOTkHKlOwLu8SPF
2IwqaFPzKBWXQczhgZTbtsWM0itBn5cB0Cws+dTJc5/24qYR2kS/6iR+E8iSdrSD
iBGh0j8TH+wbyXAo5+LvvzKNxrRjLPchXDcWosyKXwbkCRPPBW2bfN7JmkFXAHX9
F6ZDuWoJOI85YFEtkHoD0rIarbknadw476PD31ezx0f1QbRN4BK+zG+YXe1TcIfA
gHeL63gIyRwaoDq3n70/yF5o4xJ2bsmm8vT8hHoEdl5CYaO7Da9AKl94WMumH4g2
dmfzzXGYK6UTDY6xIzwTvTmFVRQeRqIAHX5Y/kzts+gBz3fvXO/EUP97YeN7exTh
cljU8v9d8a+/maWOlPzQfzl6pbwj7ef6ERlv5sD3JzRbLkGqslxgHAHnDw1Qt4dk
QN3dFFY4LOZm47NmySW+NTVTaqOE8hD/Zn9jaX2RhJkqDJZCkq8EGrpE2lzgjEbq
EwNVw93pnqWFEomQgemZV0wPb101N6thcS6cQrsQF1QSTRrtgi/JWe5vqkDQifor
9ED/TkEJcD2bszPO7yjnwo8Rr9Xuwdg2P20BA+CJM9In0kuaEUawKEBrs4gxIzXN
LKCWPZN5xGqnvcfjpBj1DioMiriF2icbTvWoIKPbIXsjhcV5pvS/yMwgxjFlyjQk
fZIkk9xWZ6QHHvTtdueIGU9+F+ENIv8B2JdhYDCJxLNeS0wzHg09qCSmWmdz4j/+
2WkojGqF6iiEnOAVxYjxDmfiCgsVThDdOwRjakEIF6soMy3wOd3lABo9PDNMJEt0
MayaOCM8L80bgfuJbbykrmJDYUn3ujKzzBN0SzkAY7fYTddod1ft/sPb2n1foo69
/e6PTUj5LwJ1vP0jcBWIPJGH4Wtq9EBm57QmVKGVf/jTDKhvqkr7ItW33ebAHILx
we8p/De7GN+ZHP2z65+tSDcb+1KFFiQBYJ1aJSRbMHuvgPEF7sRDdL3ODiMInx+b
zzmlb5qbPTdH7AbL5yF+umPgtpW/2sQgUJ4k8B0QbcsjKI5lzQbvfXGC787TJ5h/
DUgfmQg8RMgNNeRdXnsxb6ju7DB3w9tSYtWMG6gN4n4B4loKp6bqGyfEXUnWD+hE
NBJGxSk1M9W6dFf99c2/UZvwDMJ6DK6M3Eqkp5l0fz1B9c6jMkY+L+Wo70pbhyiI
aq9FEdbFm80gxmnTD1Zd5ArEhoWN2FXasOU0L4SU6BbuR+KDuGCi6uMtghoTqqeg
26uhi2OjsGEPLpuuZ2RAce5/SRbEYFHy782LmgOJfdkGCLMt55rvKOCfl60BReA7
lR+L9sFHW26aeh98G+EfJmh4xSSyi6n8uuDf+UX+8KD4pxq1NRyLHr+GsoOhGUi0
vSns0jWP6fYyXv2FzfjZf5crjyuAZ2+ndfqxaLa2DdULOI0dG+HWKC0rarY+Fm5s
nIiiCVZ5Udg6P6O4P2zKC3mC9qQhNCMp5iibGYwTELHgklzcq42QF6knEarP3NUy
tkJgY+zWh906Vth7bz5Dxhdk6OEzQ+zuxmRYfGKnqV9i7E44x7CPa/hPISR77hH8
qWrHSXUUqDG3lJF64uld9LFjNV/5Q9MqmRtZn9NNbfgdU1eShdfbf8LrEKT8PYzy
Jq1a/QfwipH+cNwzTCLAmq3FYCuOPJMMRW/YI2fQsZxUXxBLwuqrSxgl9w1Pe2vS
G9IHThAEayt785dyExEu9Ej0dew2bjmhJQz4k2wav5nH1/RCekgL+5Yb20JhsgkP
ffrGbl/iy3Br1/Jhta5sdmA8Y4PnWXEB4t1Ic6vuwyrY+4Gy2rj6fR/W8S3KQpPD
eenkm8DB3to05HrK+m4U0paHDSSR79/cYrthwWNhkCr6yovIDkk4ncOcpI0JQ2Pi
ymSlvurTCGExGCaUFMFE7hKx9adXhhToDe9zGGTl/9o51CBLNXkTnvC1GWcP2SWs
iAtW786w80hdKa08qkoyV7fTxXiDiI8PRZksZjpYaFdqy1sT/tRNfqNh82wpRZEM
czuUHEBY+sYhYU5VnA7xWuSKU9/em7pIUX4cxDO0E4AG9Lwr7wkVT42LDw5L523J
ixrH43GM0EWjIL6KIvN+ei5r/jsby43z05xHGhgXMOAmmeEzA7B4a7iK4Vpzntjv
6YtZmsoryH1oYHGBjPLOP8Bt4ztriNqhDQGHAl6gll+qH1gRaKT6BPpbXYoflUC9
nw5PM7DnK7SPWTFIwj9zH6iDKNK0qbHc4v9hjf5VNVKxwpqhH3I7rnssFTi/6b9r
thMoWgtTib67N2QUAqTjujdjMsQ4N+RWqzxSyxmm7AkcqIrT61ZiiwNgU0THE0yi
TPFAZ0RmMYFUe3Ox8m5NSk80HXBvuye928xRktubZbotvrYxBoeh4VZTA9iVOcXN
Q0zkB73seLLMN0bUVTXaoRfaKoDiv04yNTQ/bzfrazu6kIBjBXstJWQmheOYhMTW
bag/ux9HjeBnisXFel8HGYlbOhzKiHk9NIPNSRPDRZFnj1I6z7DJRL93nnA4xVtb
15wUvNamWr2zPTp87yJQfoHqA/5HGThCAMYJw0hiX6mbgEErHlT82kfPuTSGqvNm
C0H8NDLs1lCeuz14U5mJmJok/K5yHYRDPqTmPjTXgm+T65SYg1OyNRjNLgF36JT7
poYd9TjXUrxh4LtF1ImHyoNsePulY6y8SNntZUbt4LYPhEYf9L39Vx6ti+BofS2S
h4uqzpLgsX4zGcyhj/eELrucyKmsAlifpGF4qmYJQ3r/kNValEMKvi5O+zz3nsz6
niF8pgATTQioi7vuTPL2vq2xAY4Hn5r63nMijGeNL1SuhRe7LdON5axUd/cq+XRF
c+ZNjaeaEGiVyu2JEDXa9konLiTXA4MxCyCDce94+eg8pyi8cot6c0NK1W3ASyNV
FAsUf0bFbKIIkuCn2JmUORdV76xSXhpgMxqyosNnC0t5Jt4rwx/Yqx5OMA38xJKp
wHuglAXcOqSZ31pPs+xqU/tQ6YmIqRWoUi9hRH96Xb3q/lXKku5kg7zEOHAYKyAc
z9FzpFRQ2ksZv1bf+5KNhjCTKos52yvF+LIxZ80y19gBqbPYrkj/ptI3EuWWbDWI
5siK2ULz2fr+1ZW+tXS5c8nnSWwts0MQhSsPfC2xMZ8gbEaRvdi0d6XZIXGwQLCR
TANvHmzid5OM7YDGx/my4FU6IkJqz2AVCJgU43PCM15JOeNykDp2zvyDas49lpJd
CIzEyj66AS4HnO24xatRrxY6V2rLMg0GqQNTtmW6hdM7M1B9dVX2YRvtoPCyjm63
IZw0APRq+XsxOvogotQif0jWBNS2YthVw50rlzPw51BCgW2tWWIn+gkJ7Fs+fQ22
dmT87ekFu0oY7o0vw1Xa67gdDUsQf3NrHWsW3jSQ2IwXlVlZQzb50Vt5gEO+Yko0
ww5t2lEHwkbvjybqK6U8pDivefo2ffm+vYlXWazA4YtGv/Deg2knYOZY3SeyMXib
JsdJnj2z30LXihwi8Ozl+CtKsOWORAzfzqv7GdS8juNLOpOtnPgTs1yGJRnbCLfo
TcoYBdgbxwVb25cYuceoalTI3gcarUOZHsI1UklE9emIKw+zp7d0CWcmOOVDAxTr
k7Nqt47CkUbFGwExvAkOEk+qtUBOv88TCoX1cvNXI0b/kcRkOKYo7bSqA3WQ6Mx6
eGv+Qp6J9um9Q4UAhDBss/tgeH6ip+Kz4ZN8s3u4HpRfJTbtL6nj5c/L0qJb1JTM
RaCrI/3dH/6xBA79k5HdIw==
//pragma protect end_data_block
//pragma protect digest_block
mLUmyvG+NYoTOyFSd2/4eUNMqm4=
//pragma protect end_digest_block
//pragma protect end_protected
endpackage


