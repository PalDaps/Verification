
  `include "ovm_ahb_if_wrapper.sv"
  `include "ovm_ahb_tran_item.sv"
  `include "ovm_ahb_master_driver.sv"
  `include "ovm_ahb_master_sequencer.sv"
  `include "ovm_ahb_seq_lib.sv"
  `include "ovm_ahb_monitor.sv"
  `include "ovm_ahb_agent.sv"