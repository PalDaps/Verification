// $Id: ovm_in_order_comparator.svh,v 1.11 2009/05/12 21:02:29 redelman Exp $
//------------------------------------------------------------------------------
//   Copyright 2007-2009 Mentor Graphics Corporation
//   Copyright 2007-2009 Cadence Design Systems, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
//
// CLASS: ovm_in_order_comparator #(T,comp_type,convert,pair_type)
//
// Compares two streams of data objects of type T, a parameter to this class.
// These transactions may either be classes or built-in types. To be
// successfully compared, the two streams of data must be in the same order.
// Apart from that, there are no assumptions made about the relative timing of
// the two streams of data.
//
// Type parameters
//
//   T       - Specifies the type of transactions to be compared.
//
//   comp    - The type of the comparator to be used to compare the two
//             transaction streams.
//
//   convert - A policy class to allow convert2string() to be called on the
//             transactions being compared. If T is an extension of
//             ovm_transaction, then it uses T::convert2string(). If T is a
//             built-in type, then the policy provides a convert2string()
//             method for the comparator to call. 
//
//  pair_type - A policy class to allow pairs of transactions to be handled as
//             a single ovm_transaction type.
//
// Built in types (such as ints, bits, logic, and structs) can be compared using
// the default values for comp_type, convert, and pair_type. For convenience,
// you can use the subtype, <ovm_in_order_builtin_comparator #(T)> for built-in
// types.
//
// When T is a class, T must implement comp and convert2string, and you must
// specify class-based policy classes for comp_type, convert, and pair_type.
// In most cases, you can use the convenient subtype,
// ovm_in_order_class_comparator #(T).
//
// Comparisons are commutative, meaning it does not matter which data stream is
// connected to which export, before_export or after_export.
//
// Comparisons are done in order and as soon as a transaction is received from
// both streams. Internal fifos are used to buffer incoming transactions on one
// stream until a transaction to compare arrives on the other stream.
//
//------------------------------------------------------------------------------

class ovm_in_order_comparator 
  #( type T = int ,
     type comp_type = ovm_built_in_comp #( T ) ,
     type convert = ovm_built_in_converter #( T ) , 
     type pair_type = ovm_built_in_pair #( T ) )
    extends ovm_component;

  typedef ovm_in_order_comparator #(T,comp_type,convert,pair_type) this_type;
  `ovm_component_param_utils(this_type)

  const static string type_name = 
    "ovm_in_order_comparator #(T,comp_type,convert,pair_type)";

  // Port: before_export
  //
  // The export to which one stream of data is written. The port must be
  // connected to an analysis port that will provide such data. 

  ovm_analysis_export #(T) before_export;


  // Port: after_export
  //
  // The export to which the other stream of data is written. The port must be
  // connected to an analysis port that will provide such data. 

  ovm_analysis_export #(T) after_export;


  // Port: pair_ap
  //
  // The comparator sends out pairs of transactions across this analysis port.
  // Both matched and unmatched pairs are published via a pair_type objects.
  // Any connected analysis export(s) will receive these transaction pairs.

  ovm_analysis_port   #(pair_type) pair_ap;
  
  local tlm_analysis_fifo #(T) m_before_fifo;
  local tlm_analysis_fifo #(T) m_after_fifo;

  int m_matches, m_mismatches;

  function new(string name, ovm_component parent);

    super.new(name, parent);

    before_export = new("before_export", this);
    after_export  = new("after_export", this);
    pair_ap       = new("pair_ap", this);

    m_before_fifo = new("before", this);
    m_after_fifo  = new("after", this);
    m_matches = 0;
    m_mismatches = 0;

  endfunction
  
  virtual function string get_type_name();
    return type_name;
  endfunction

  virtual function void connect();
    before_export.connect(m_before_fifo.analysis_export);
    after_export.connect(m_after_fifo.analysis_export);
  endfunction


  // Task- run
  //
  // Internal method.
  //
  // Takes pairs of before and after transactions and compares them. 
  // Status information is updated according to the results of the comparison.
  // Each pair is published to the pair_ap analysis port.

  virtual task run();
 
    pair_type pair;
    T b;
    T a;
  
    string s;
   
    forever begin
      
      m_before_fifo.get(b);
      m_after_fifo.get(a);
      
      if(!comp_type::comp(b, a)) begin

        $sformat(s, "%s differs from %s", convert::convert2string(a),
                                          convert::convert2string(b));

        ovm_report_warning("Comparator Mismatch", s);

        m_mismatches++;

      end
      else begin
        s = convert::convert2string(b);
        if(ovm_report_enabled(OVM_MEDIUM))
          ovm_report_info("Comparator Match", s, OVM_MEDIUM);
        m_matches++;
      end

      // we make the assumption here that a transaction "sent for
      // analysis" is safe from being edited by another process.
      // Hence, it is safe not to clone a and b.
      
      pair = new(a, b);
      pair_ap.write(pair);
    end
  
  endtask


  // Function: flush
  //
  // This method sets m_matches and m_mismatches back to zero. The
  // <tlm_fifo #(T)::flush> takes care of flushing the FIFOs.

  virtual function void flush();
    m_matches = 0;
    m_mismatches = 0;
  endfunction
  
endclass


//------------------------------------------------------------------------------
//
// CLASS: in_order_built_in_comparator #(T)
//
// This class uses the ovm_built_in_* comparison, converter, and pair classes.
// Use this class for built-in types (int, bit, string, etc.)
//
//------------------------------------------------------------------------------

class ovm_in_order_built_in_comparator #(type T=int)
  extends ovm_in_order_comparator #(T);

  typedef ovm_in_order_built_in_comparator #(T) this_type;
  `ovm_component_param_utils(this_type)

  const static string type_name = "ovm_in_order_built_in_comparator #(T)";

  function new(string name, ovm_component parent);
    super.new(name, parent);
  endfunction
  
  virtual function string get_type_name ();
    return type_name;
  endfunction

endclass


//------------------------------------------------------------------------------
//
// CLASS: in_order_class_comparator #(T)
//
// This class uses the ovm_class_* comparison, converter, and pair classes.
// Use this class for comparing user-defined objects of type T, which must
// provide implementations of comp and convert2string.
//
//------------------------------------------------------------------------------

class ovm_in_order_class_comparator #( type T = int )
  extends ovm_in_order_comparator #( T , 
                                     ovm_class_comp #( T ) , 
                                     ovm_class_converter #( T ) , 
                                     ovm_class_pair #( T, T ) );

  typedef ovm_in_order_class_comparator #(T) this_type;
  `ovm_component_param_utils(this_type)

  const static string type_name = "ovm_in_order_class_comparator #(T)";

  function new( string name  , ovm_component parent);
    super.new( name, parent );
  endfunction
  
  virtual function string get_type_name ();
    return type_name;
  endfunction

endclass
