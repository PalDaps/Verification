//--------------------------- IP_CORE_LABS-------------------------------------//
//                        SPI_TX example project                               //
//                        file -  test_files.sv                                //
//                        harness file list                                    //
//                        author -  fputrya                                    //
//-----------------------------------------------------------------------------//

import ovm_pkg::*;

`include "ovm_macros.svh"

`include "ovm_ahb_vc_files.sv"
`include "ovm_spi_vc_files.sv"
`include "ovm_design_spec_files.sv"
`include "harness.sv"