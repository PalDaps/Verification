//--------------------------- IP_CORE_LABS-------------------------------------//
//                        SPI_TX example project                               //
//                        file -  ovm_design_spec.sv                           //
//                        design specific stuff filelist                       //
//                        author -  fputrya                                    //
//-----------------------------------------------------------------------------//

`ifndef OVM_DESIGN_SPEC
`define OVM_DESIGN_SPEC

  import ovm_pkg::*;
  `include "ovm_macros.svh"
  `include "ovm_design_spec_class_files.sv"

`endif