`ifndef OVM_SPI_VC_PKG
`define OVM_SPI_VC_PKG

`include "spi_if.sv"

package ovm_spi_vc_pkg;

   import ovm_pkg::*;
  `include "ovm_macros.svh"

  `include "ovm_spi_vc_class_files.sv"

endpackage

`endif