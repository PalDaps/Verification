//--------------------------- IP_CORE_LABS-------------------------------------//
//                        SPI_TX example project                               //
//                        file -  ovm_ahb_vc_files.sv                          //
//                        ahb verification component filelist                  //
//                        author -  fputrya                                    //
//-----------------------------------------------------------------------------//

`ifndef OVM_AHB_VC
`define OVM_AHB_VC

  `include "ahb_if.sv"

   import ovm_pkg::*;
  `include "ovm_macros.svh"
  `include "ovm_ahb_vc_class_files.sv"

`endif