//--------------------------- IP_CORE_LABS-------------------------------------//
//                        SPI_TX example project                               //
//                        file -  ovm_spi_vc_files.sv                          //
//                        spi agent file list                                  //
//                        author -  fputrya                                    //
//-----------------------------------------------------------------------------//

`ifndef OVM_SPI_VC
`define OVM_SPI_VC

  `include "spi_if.sv"

   import ovm_pkg::*;
  `include "ovm_macros.svh"

  `include "ovm_spi_vc_class_files.sv"

`endif