//----------------------------------------------------------------------
//   Copyright 2007-2009 Mentor Graphics Corporation
//   Copyright 2007-2009 Cadence Design Systems, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------
// This file undefs all macros that are defined by the OVM library. This can
// be used to load ovm into multiple scopes using a single compilation.

`undef ANSI_BG_BLACK
`undef ANSI_BG_BLUE
`undef ANSI_BG_CYAN
`undef ANSI_BG_GREEN
`undef ANSI_BG_MAGENTA
`undef ANSI_BG_RED
`undef ANSI_BG_WHITE
`undef ANSI_BG_YELLOW
`undef ANSI_BOLD
`undef ANSI_BRIGHT
`undef ANSI_DIM
`undef ANSI_FG_BLACK
`undef ANSI_FG_BLUE
`undef ANSI_FG_CYAN
`undef ANSI_FG_GREEN
`undef ANSI_FG_MAGENTA
`undef ANSI_FG_RED
`undef ANSI_FG_WHITE
`undef ANSI_FG_YELLOW
`undef ANSI_RESET
`undef ANSI_REVERSE
`undef ANSI_UNDERSCORE
`undef AVM_PKG_SV
`undef AVM_compatibility_SVH
`undef BACKWARD_COMPAT_MACROS_SVH
`undef BASE_COMPATIBILITY_SVH
`undef BLOCKING_GET_IMP
`undef BLOCKING_GET_IMP_SFX
`undef BLOCKING_PEEK_IMP
`undef BLOCKING_PEEK_IMP_SFX
`undef BLOCKING_PUT_IMP
`undef BLOCKING_PUT_IMP_SFX
`undef BLOCKING_TRANSPORT_IMP
`undef BLOCKING_TRANSPORT_IMP_SFX
`undef CDNS_RECORDING_SVH
`undef CDNS_TCL_INTERFACE_SVH
`undef COMPATIBILITY_SVH
`undef DODEEPCOPY
`undef DOREFERENCECOPY
`undef DOSHALLOWCOPY
`undef DUT_ERROR
`undef FUNCTION_ERROR
`undef MESSAGE
`undef NONBLOCKING_GET_IMP
`undef NONBLOCKING_GET_IMP_SFX
`undef NONBLOCKING_PEEK_IMP
`undef NONBLOCKING_PEEK_IMP_SFX
`undef NONBLOCKING_PUT_IMP
`undef NONBLOCKING_PUT_IMP_SFX
`undef NONBLOCKING_TRANSPORT_IMP
`undef NONBLOCKING_TRANSPORT_IMP_SFX
`undef OVM_AGENT_SVH
`undef OVM_APPLY_CONFIG_SETTING
`undef OVM_USE_SFORMATF
`undef OVM_BASE_ONLY
`undef OVM_BASE_PKG_SV
`undef OVM_BASE_SVH
`undef OVM_COMPARE_FAILED
`undef OVM_COMPONENT_SVH
`undef OVM_CONNECTOR_BASE_SVH
`undef OVM_DRIVER_SVH
`undef OVM_ENUM
`undef OVM_ENV_SVH
`undef OVM_EVENT_SVH
`undef OVM_EXTERN_REPORT_SERVER_SVH
`undef OVM_FACTORY_SVH
`undef OVM_FIELD_DATA
`undef OVM_FIELD_DATA_AA_generic
`undef OVM_FIELD_DATA_AA_int_key
`undef OVM_FIELD_DATA_AA_int_string
`undef OVM_FIELD_DATA_AA_object_int
`undef OVM_FIELD_DATA_AA_object_string
`undef OVM_FIELD_DATA_AA_string_string
`undef OVM_FIELD_DATA_ARRAY
`undef OVM_FIELD_DATA_ARRAY_OBJECT
`undef OVM_FIELD_DATA_ARRAY_STRING
`undef OVM_FIELD_DATA_EVENT
`undef OVM_FIELD_DATA_OBJECT
`undef OVM_FIELD_DATA_SARRAY
`undef OVM_FIELD_DATA_STRING
`undef OVM_FIELD_ENUM
`undef OVM_FIELD_SET
`undef OVM_FIELD_SET_AA_INT_TYPE
`undef OVM_FIELD_SET_AA_OBJECT_TYPE
`undef OVM_FIELD_SET_AA_TYPE
`undef OVM_FIELD_SET_ARRAY_OBJECT
`undef OVM_FIELD_SET_ARRAY_OBJECT_TYPE
`undef OVM_FIELD_SET_ARRAY_TYPE
`undef OVM_FIELD_SET_EVENT
`undef OVM_FIELD_SET_OBJECT
`undef OVM_FIELD_SET_QUEUE_OBJECT
`undef OVM_FIELD_SET_QUEUE_OBJECT_TYPE
`undef OVM_FIELD_SET_QUEUE_TYPE
`undef OVM_FIELD_SET_STRING
`undef OVM_LINE_WIDTH
`undef OVM_LOCAL_SCOPE_STACK
`undef OVM_MACROS_SVH
`undef OVM_METH_DEFINES_SVH
`undef OVM_METH_SVH
`undef OVM_MISC_SVH
`undef OVM_MONITOR_SVH
`undef OVM_NUM_LINES
`undef OVM_OBJECT_DEFINES_SVH
`undef OVM_OBJECT_GLOBALS_SVH
`undef OVM_OBJECT_SVH
`undef OVM_PACKER_SVH
`undef OVM_PAIR_SVH
`undef OVM_PHASES_SVH
`undef OVM_PHASE_EVENT_CB_TASK
`undef OVM_PKG_SV
`undef OVM_POLICIES_SVH
`undef OVM_PRINTER_DEFINES_SVH
`undef OVM_PRINTER_SVH
`undef OVM_RECORD_INTERFACE
`undef OVM_REGISTRY_SVH
`undef OVM_REPORT_CLIENT_SVH
`undef OVM_REPORT_DEFINES_SVH
`undef OVM_REPORT_GLOBAL_SVH
`undef OVM_REPORT_HANDLER_SVH
`undef OVM_REPORT_SERVER_SVH
`undef OVM_REQ_RSP_DRIVER_SVH
`undef OVM_REQ_RSP_SEQUENCE_SVH
`undef OVM_SCOREBOARD_SVH
`undef OVM_SEQUENCER_BASE_SVH
`undef OVM_SEQUENCER_SVH
`undef OVM_SEQUENCE_BUILTIN_SVH
`undef OVM_SEQUENCE_ITEM_SVH
`undef OVM_SEQUENCE_SVH
`undef OVM_SVH
`undef OVM_TEST_SVH
`undef OVM_THREADED_COMPONENT_SVH
`undef OVM_TRANSACTION_SVH
`undef OVM_URM_MESSAGE_DEFINES_SVH
`undef OVM_URM_MESSAGE_SVH
`undef OVM_VERSION_SVH
`undef OVM_VIRTUAL_SEQUENCER_SVH
`undef RESIZE_QUEUE_COPY
`undef RESIZE_QUEUE_NOCOPY
`undef RESIZE_QUEUE_OBJECT_COPY
`undef RESIZE_QUEUE_OBJECT_NOCOPY
`undef TASK_ERROR
`undef TLM_ANALYSIS_MASK
`undef TLM_BLOCKING_GET_MASK
`undef TLM_BLOCKING_GET_PEEK_MASK
`undef TLM_BLOCKING_MASTER_MASK
`undef TLM_BLOCKING_PEEK_MASK
`undef TLM_BLOCKING_PUT_MASK
`undef TLM_BLOCKING_SLAVE_MASK
`undef TLM_BLOCKING_TRANSPORT_MASK
`undef TLM_FIFO_FUNCTION_ERROR
`undef TLM_FIFO_TASK_ERROR
`undef TLM_GET_MASK
`undef TLM_GET_PEEK_MASK
`undef TLM_MASTER_MASK
`undef TLM_NONBLOCKING_GET_MASK
`undef TLM_NONBLOCKING_GET_PEEK_MASK
`undef TLM_NONBLOCKING_PEEK_MASK
`undef TLM_NONBLOCKING_PUT_MASK
`undef TLM_NONBLOCKING_SLAVE_MASK
`undef TLM_NONBLOCKING_TRANSPORT_MASK
`undef TLM_PEEK_MASK
`undef TLM_PUT_MASK
`undef TLM_SLAVE_MASK
`undef TLM_TRANSPORT_MASK
`undef URM_GLOBALS
`undef URM_METH_COMPATIBILITY_SVH
`undef URM_SVH
`undef URM_TYPE_COMPATIBILITY_SVH
`undef abstract_avm_to_ovm_component
`undef avm_to_ovm_bidi
`undef avm_to_ovm_component
`undef avm_to_ovm_policy
`undef avm_to_ovm_uni
`undef cdns_ovm_major_rev
`undef cdns_ovm_minor_rev
`undef cdns_ovm_name
`undef cdns_ovm_sub_rev
`undef const
`undef dut_error
`undef extern
`undef local
`undef message
`undef ovm_analysis_imp_decl
`undef ovm_blocking_get_imp_decl
`undef ovm_blocking_get_peek_imp_decl
`undef ovm_blocking_master_imp_decl
`undef ovm_blocking_peek_imp_decl
`undef ovm_blocking_put_imp_decl
`undef ovm_blocking_slave_imp_decl
`undef ovm_blocking_transport_imp_decl
`undef ovm_factory_override_func
`undef ovm_component_factory_create_func
`undef ovm_component_new_func
`undef ovm_component_registry
`undef ovm_component_registry_param
`undef ovm_component_registry_internal
`undef ovm_component_utils
`undef ovm_component_utils_begin
`undef ovm_component_utils_end
`undef ovm_create
`undef ovm_create_seq
`undef ovm_declare_sequence_lib
`undef ovm_do
`undef ovm_do_seq
`undef ovm_do_seq_with
`undef ovm_do_with
`undef ovm_end_package
`undef ovm_error
`undef ovm_fatal
`undef ovm_field_aa_int_byte
`undef ovm_field_aa_int_byte_unsigned
`undef ovm_field_aa_int_int
`undef ovm_field_aa_int_int_unsigned
`undef ovm_field_aa_int_integer
`undef ovm_field_aa_int_integer_unsigned
`undef ovm_field_aa_int_key
`undef ovm_field_aa_int_longint
`undef ovm_field_aa_int_longint_unsigned
`undef ovm_field_aa_int_shortint
`undef ovm_field_aa_int_shortint_unsigned
`undef ovm_field_aa_int_string
`undef ovm_field_aa_object_int
`undef ovm_field_aa_object_string
`undef ovm_field_aa_string_int
`undef ovm_field_aa_string_string
`undef ovm_field_array_int
`undef ovm_field_array_object
`undef ovm_field_array_string
`undef ovm_field_enum
`undef ovm_field_event
`undef ovm_field_int
`undef ovm_field_object
`undef ovm_field_queue_int
`undef ovm_field_queue_object
`undef ovm_field_queue_string
`undef ovm_field_sarray_int
`undef ovm_field_string
`undef ovm_field_utils
`undef ovm_field_utils_begin
`undef ovm_field_utils_end
`undef ovm_file
`undef ovm_get_imp_decl
`undef ovm_get_peek_imp_decl
`undef ovm_get_type_name_func
`undef ovm_global_reporter
`undef ovm_global_urm_report_server
`undef ovm_info
`undef ovm_line
`undef ovm_master_imp_decl
`undef ovm_msg_detail
`undef ovm_named_object_create_func
`undef ovm_named_object_factory_create_func
`undef ovm_named_object_new_func
`undef ovm_new_func
`undef ovm_new_func_data
`undef ovm_non_blocking_transport_imp_decl
`undef ovm_nonblocking_get_imp_decl
`undef ovm_nonblocking_get_peek_imp_decl
`undef ovm_nonblocking_master_imp_decl
`undef ovm_nonblocking_peek_imp_decl
`undef ovm_nonblocking_put_imp_decl
`undef ovm_nonblocking_slave_imp_decl
`undef ovm_object_create_func
`undef ovm_object_factory_create_func
`undef ovm_object_new_func
`undef ovm_object_registry
`undef ovm_object_registry_param
`undef ovm_object_registry_internal
`undef ovm_object_utils
`undef ovm_object_utils_begin
`undef ovm_object_utils_end
`undef ovm_package
`undef ovm_packages
`undef ovm_peek_imp_decl
`undef ovm_phase_func_decl
`undef ovm_phase_task_decl
`undef ovm_print_aa_int_key4
`undef ovm_print_aa_int_object
`undef ovm_print_aa_int_object3
`undef ovm_print_aa_string_int
`undef ovm_print_aa_string_int3
`undef ovm_print_aa_string_object
`undef ovm_print_aa_string_object3
`undef ovm_print_aa_string_string
`undef ovm_print_aa_string_string2
`undef ovm_print_array_int
`undef ovm_print_array_int3
`undef ovm_print_array_object
`undef ovm_print_array_object3
`undef ovm_print_array_string
`undef ovm_print_array_string2
`undef ovm_print_int
`undef ovm_print_int3
`undef ovm_print_msg_enum
`undef ovm_print_object
`undef ovm_print_object2
`undef ovm_print_object_qda4
`undef ovm_print_object_queue
`undef ovm_print_object_queue3
`undef ovm_print_qda_int4
`undef ovm_print_queue_int
`undef ovm_print_queue_int3
`undef ovm_print_string
`undef ovm_print_string2
`undef ovm_print_string_qda3
`undef ovm_print_string_queue
`undef ovm_print_string_queue2
`undef ovm_put_imp_decl
`undef ovm_rand_send
`undef ovm_rand_send_with
`undef ovm_record_any_object
`undef ovm_record_array_int
`undef ovm_record_array_object
`undef ovm_record_array_string
`undef ovm_record_int
`undef ovm_record_object
`undef ovm_record_string
`undef ovm_register_self_func
`undef ovm_register_sequence
`undef ovm_send
`undef ovm_sequence_library_package
`undef ovm_sequence_utils
`undef ovm_sequence_utils_begin
`undef ovm_sequence_utils_end
`undef ovm_sequencer_utils
`undef ovm_sequencer_utils_begin
`undef ovm_sequencer_utils_end
`undef ovm_set_flags
`undef ovm_slave_imp_decl
`undef ovm_transport_imp_decl
`undef ovm_update_sequence_lib
`undef ovm_update_sequence_lib_and_item
`undef ovm_urm_message
`undef ovm_urm_report_server
`undef ovm_urm_reporter
`undef ovm_urm_tmp_str
`undef ovm_warning
`undef print_integral_field
`undef ref
`undef static_dut_error
`undef static_message
`undef tlm_export_compat_new_func
`undef tlm_port_compat_new_func
`undef urm_code_debug
`undef urm_component_factory_create_func
`undef urm_data_debug
`undef urm_debug
`undef urm_error
`undef urm_error_id
`undef urm_fatal
`undef urm_fatal_id
`undef urm_field_aa_int_byte
`undef urm_field_aa_int_byte_unsigned
`undef urm_field_aa_int_int
`undef urm_field_aa_int_int_unsigned
`undef urm_field_aa_int_integer
`undef urm_field_aa_int_integer_unsigned
`undef urm_field_aa_int_key
`undef urm_field_aa_int_longint
`undef urm_field_aa_int_longint_unsigned
`undef urm_field_aa_int_shortint
`undef urm_field_aa_int_shortint_unsigned
`undef urm_field_aa_int_string
`undef urm_field_aa_object_int
`undef urm_field_aa_object_string
`undef urm_field_aa_string_string
`undef urm_field_array_int
`undef urm_field_array_object
`undef urm_field_array_string
`undef urm_field_event
`undef urm_field_int
`undef urm_field_object
`undef urm_field_queue_int
`undef urm_field_queue_object
`undef urm_field_queue_string
`undef urm_field_string
`undef urm_field_utils
`undef urm_field_utils_begin
`undef urm_field_utils_end
`undef urm_file
`undef urm_flow_debug
`undef urm_info
`undef urm_info0
`undef urm_info1
`undef urm_info2
`undef urm_info3
`undef urm_info4
`undef urm_info_id
`undef urm_line
`undef urm_msg_detail
`undef urm_msg_imp
`undef urm_object_utils
`undef urm_object_utils_begin
`undef urm_object_utils_end
`undef urm_pkg_msg_imp
`undef urm_static_code_debug
`undef urm_static_data_debug
`undef urm_static_debug
`undef urm_static_error
`undef urm_static_error_id
`undef urm_static_fatal
`undef urm_static_fatal_id
`undef urm_static_flow_debug
`undef urm_static_info
`undef urm_static_info0
`undef urm_static_info1
`undef urm_static_info2
`undef urm_static_info3
`undef urm_static_info4
`undef urm_static_info_id
`undef urm_static_msg_detail
`undef urm_static_warning
`undef urm_static_warning_id
`undef urm_unit_base_utils
`undef urm_unit_base_utils_begin
`undef urm_unit_base_utils_end
`undef urm_unit_utils
`undef urm_unit_utils_begin
`undef urm_unit_utils_end
`undef urm_unit_wrapper_derived_class
`undef urm_warning
`undef urm_warning_id
