//----------------------------------------------------------------------
//   Copyright 2007-2009 Cadence Design Systems, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------

`ifndef CDNS_ADDITIONS_SVH
`define CDNS_ADDITIONS_SVH

`ifdef INCA
  `include "cdns_additions/cdns_recording.svh"
  `include "cdns_additions/cdns_tcl_interface.svh"
`endif

  `include "cdns_additions/ovm_mb_utils.sv"

`endif // CDNS_ADDITIONS_SVH
